
library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic
	(
		ADDR_WIDTH : integer := 15 -- Specify your actual ROM size to save LEs and unnecessary block RAM usage.
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture rtl of controller_rom1 is

	signal addr1 : integer range 0 to 2**ADDR_WIDTH-1;

	--  build up 2D array to hold the memory
	type word_t is array (0 to 3) of std_logic_vector(7 downto 0);
	type ram_t is array (0 to 2 ** ADDR_WIDTH - 1) of word_t;

	signal ram : ram_t:=
	(

     0 => (x"04",x"87",x"da",x"01"),
     1 => (x"58",x"0e",x"87",x"dd"),
     2 => (x"0e",x"5a",x"59",x"5e"),
     3 => (x"00",x"00",x"29",x"27"),
     4 => (x"4a",x"26",x"0f",x"00"),
     5 => (x"48",x"26",x"49",x"26"),
     6 => (x"08",x"26",x"80",x"ff"),
     7 => (x"00",x"2d",x"27",x"4f"),
     8 => (x"27",x"4f",x"00",x"00"),
     9 => (x"00",x"00",x"00",x"2a"),
    10 => (x"fd",x"00",x"4f",x"4f"),
    11 => (x"fc",x"f7",x"c4",x"87"),
    12 => (x"86",x"c0",x"c5",x"4e"),
    13 => (x"49",x"fc",x"f7",x"c4"),
    14 => (x"48",x"c4",x"fe",x"c3"),
    15 => (x"40",x"40",x"c0",x"89"),
    16 => (x"89",x"d0",x"40",x"40"),
    17 => (x"c1",x"87",x"f6",x"03"),
    18 => (x"00",x"87",x"fa",x"f0"),
    19 => (x"1e",x"87",x"fc",x"98"),
    20 => (x"48",x"12",x"1e",x"72"),
    21 => (x"87",x"c4",x"02",x"11"),
    22 => (x"87",x"f6",x"02",x"88"),
    23 => (x"4f",x"26",x"4a",x"26"),
    24 => (x"73",x"1e",x"72",x"1e"),
    25 => (x"11",x"48",x"12",x"1e"),
    26 => (x"4b",x"87",x"ca",x"02"),
    27 => (x"9b",x"98",x"df",x"c3"),
    28 => (x"f0",x"02",x"88",x"73"),
    29 => (x"26",x"4b",x"26",x"87"),
    30 => (x"1e",x"4f",x"26",x"4a"),
    31 => (x"1e",x"72",x"1e",x"73"),
    32 => (x"ca",x"04",x"8b",x"c1"),
    33 => (x"11",x"48",x"12",x"87"),
    34 => (x"88",x"87",x"c4",x"02"),
    35 => (x"26",x"87",x"f1",x"02"),
    36 => (x"26",x"4b",x"26",x"4a"),
    37 => (x"1e",x"74",x"1e",x"4f"),
    38 => (x"1e",x"72",x"1e",x"73"),
    39 => (x"d0",x"04",x"8b",x"c1"),
    40 => (x"11",x"48",x"12",x"87"),
    41 => (x"4c",x"87",x"ca",x"02"),
    42 => (x"9c",x"98",x"df",x"c3"),
    43 => (x"eb",x"02",x"88",x"74"),
    44 => (x"26",x"4a",x"26",x"87"),
    45 => (x"26",x"4c",x"26",x"4b"),
    46 => (x"48",x"73",x"1e",x"4f"),
    47 => (x"02",x"a9",x"73",x"81"),
    48 => (x"53",x"12",x"87",x"c5"),
    49 => (x"26",x"87",x"f6",x"05"),
    50 => (x"48",x"73",x"1e",x"4f"),
    51 => (x"05",x"a9",x"73",x"81"),
    52 => (x"87",x"f9",x"53",x"72"),
    53 => (x"5e",x"0e",x"4f",x"26"),
    54 => (x"0e",x"5d",x"5c",x"5b"),
    55 => (x"4d",x"71",x"86",x"f4"),
    56 => (x"c0",x"48",x"a6",x"c4"),
    57 => (x"4b",x"66",x"dc",x"78"),
    58 => (x"c0",x"48",x"a6",x"c8"),
    59 => (x"7e",x"97",x"15",x"78"),
    60 => (x"c0",x"02",x"6e",x"97"),
    61 => (x"4c",x"13",x"87",x"f0"),
    62 => (x"87",x"da",x"02",x"9c"),
    63 => (x"74",x"4a",x"6e",x"97"),
    64 => (x"05",x"aa",x"b7",x"49"),
    65 => (x"a6",x"c8",x"87",x"c9"),
    66 => (x"c0",x"78",x"c1",x"48"),
    67 => (x"13",x"87",x"c2",x"4c"),
    68 => (x"05",x"9c",x"74",x"4c"),
    69 => (x"66",x"c8",x"87",x"e6"),
    70 => (x"c4",x"87",x"cb",x"02"),
    71 => (x"80",x"c1",x"48",x"66"),
    72 => (x"fe",x"58",x"a6",x"c8"),
    73 => (x"66",x"c4",x"87",x"ff"),
    74 => (x"26",x"8e",x"f4",x"48"),
    75 => (x"26",x"4c",x"26",x"4d"),
    76 => (x"1e",x"4f",x"26",x"4b"),
    77 => (x"c1",x"c1",x"4a",x"71"),
    78 => (x"d9",x"04",x"aa",x"b7"),
    79 => (x"b7",x"c6",x"c1",x"87"),
    80 => (x"87",x"d2",x"01",x"aa"),
    81 => (x"d0",x"48",x"66",x"c4"),
    82 => (x"87",x"ca",x"05",x"a8"),
    83 => (x"f7",x"c0",x"49",x"72"),
    84 => (x"c0",x"48",x"71",x"89"),
    85 => (x"e1",x"c1",x"87",x"ec"),
    86 => (x"d8",x"04",x"aa",x"b7"),
    87 => (x"b7",x"e6",x"c1",x"87"),
    88 => (x"87",x"d1",x"01",x"aa"),
    89 => (x"d0",x"48",x"66",x"c4"),
    90 => (x"87",x"c9",x"05",x"a8"),
    91 => (x"d7",x"c1",x"49",x"72"),
    92 => (x"cd",x"48",x"71",x"89"),
    93 => (x"8a",x"f0",x"c0",x"87"),
    94 => (x"06",x"aa",x"b7",x"c9"),
    95 => (x"4a",x"ff",x"87",x"c2"),
    96 => (x"4f",x"26",x"48",x"72"),
    97 => (x"5c",x"5b",x"5e",x"0e"),
    98 => (x"86",x"f8",x"0e",x"5d"),
    99 => (x"a6",x"c4",x"7e",x"71"),
   100 => (x"4c",x"78",x"c0",x"48"),
   101 => (x"1e",x"a7",x"f9",x"c1"),
   102 => (x"fc",x"49",x"66",x"c4"),
   103 => (x"86",x"c4",x"87",x"f8"),
   104 => (x"4b",x"6e",x"49",x"70"),
   105 => (x"6b",x"97",x"83",x"71"),
   106 => (x"a9",x"ed",x"c0",x"49"),
   107 => (x"c4",x"87",x"c6",x"05"),
   108 => (x"78",x"c1",x"48",x"a6"),
   109 => (x"02",x"66",x"d8",x"83"),
   110 => (x"66",x"d8",x"87",x"c5"),
   111 => (x"97",x"0b",x"7b",x"0b"),
   112 => (x"87",x"d3",x"05",x"6b"),
   113 => (x"c7",x"02",x"66",x"c4"),
   114 => (x"c0",x"4a",x"74",x"87"),
   115 => (x"87",x"c2",x"8a",x"0a"),
   116 => (x"48",x"72",x"4a",x"74"),
   117 => (x"dc",x"87",x"ef",x"c0"),
   118 => (x"49",x"13",x"1e",x"66"),
   119 => (x"c4",x"87",x"d4",x"fd"),
   120 => (x"c0",x"4d",x"70",x"86"),
   121 => (x"d4",x"03",x"ad",x"b7"),
   122 => (x"02",x"66",x"c4",x"87"),
   123 => (x"48",x"74",x"87",x"c9"),
   124 => (x"70",x"88",x"08",x"c0"),
   125 => (x"74",x"87",x"c2",x"7e"),
   126 => (x"c9",x"48",x"6e",x"7e"),
   127 => (x"94",x"66",x"dc",x"87"),
   128 => (x"fe",x"4c",x"a4",x"75"),
   129 => (x"8e",x"f8",x"87",x"ef"),
   130 => (x"4c",x"26",x"4d",x"26"),
   131 => (x"4f",x"26",x"4b",x"26"),
   132 => (x"73",x"1e",x"00",x"20"),
   133 => (x"02",x"9a",x"72",x"1e"),
   134 => (x"c0",x"87",x"e7",x"c0"),
   135 => (x"72",x"4b",x"c1",x"48"),
   136 => (x"87",x"d1",x"06",x"a9"),
   137 => (x"c9",x"06",x"82",x"72"),
   138 => (x"72",x"83",x"73",x"87"),
   139 => (x"87",x"f4",x"01",x"a9"),
   140 => (x"b2",x"c1",x"87",x"c3"),
   141 => (x"03",x"a9",x"72",x"3a"),
   142 => (x"07",x"80",x"73",x"89"),
   143 => (x"05",x"2b",x"2a",x"c1"),
   144 => (x"4b",x"26",x"87",x"f3"),
   145 => (x"75",x"1e",x"4f",x"26"),
   146 => (x"71",x"4d",x"c4",x"1e"),
   147 => (x"ff",x"04",x"a1",x"b7"),
   148 => (x"c3",x"81",x"c1",x"b9"),
   149 => (x"b7",x"72",x"07",x"bd"),
   150 => (x"ba",x"ff",x"04",x"a2"),
   151 => (x"bd",x"c1",x"82",x"c1"),
   152 => (x"87",x"ee",x"fe",x"07"),
   153 => (x"ff",x"04",x"2d",x"c1"),
   154 => (x"07",x"80",x"c1",x"b8"),
   155 => (x"b9",x"ff",x"04",x"2d"),
   156 => (x"26",x"07",x"81",x"c1"),
   157 => (x"1e",x"4f",x"26",x"4d"),
   158 => (x"4a",x"71",x"1e",x"73"),
   159 => (x"49",x"4b",x"66",x"c8"),
   160 => (x"99",x"71",x"8b",x"c1"),
   161 => (x"12",x"87",x"cf",x"02"),
   162 => (x"08",x"d4",x"ff",x"48"),
   163 => (x"c1",x"49",x"73",x"78"),
   164 => (x"05",x"99",x"71",x"8b"),
   165 => (x"4b",x"26",x"87",x"f1"),
   166 => (x"5e",x"0e",x"4f",x"26"),
   167 => (x"71",x"0e",x"5c",x"5b"),
   168 => (x"4c",x"d4",x"ff",x"4a"),
   169 => (x"49",x"4b",x"66",x"cc"),
   170 => (x"99",x"71",x"8b",x"c1"),
   171 => (x"c3",x"87",x"ce",x"02"),
   172 => (x"52",x"6c",x"7c",x"ff"),
   173 => (x"8b",x"c1",x"49",x"73"),
   174 => (x"f2",x"05",x"99",x"71"),
   175 => (x"26",x"4c",x"26",x"87"),
   176 => (x"1e",x"4f",x"26",x"4b"),
   177 => (x"d4",x"ff",x"1e",x"73"),
   178 => (x"7b",x"ff",x"c3",x"4b"),
   179 => (x"ff",x"c3",x"4a",x"6b"),
   180 => (x"c8",x"49",x"6b",x"7b"),
   181 => (x"c3",x"b1",x"72",x"32"),
   182 => (x"4a",x"6b",x"7b",x"ff"),
   183 => (x"b2",x"71",x"31",x"c8"),
   184 => (x"6b",x"7b",x"ff",x"c3"),
   185 => (x"72",x"32",x"c8",x"49"),
   186 => (x"26",x"48",x"71",x"b1"),
   187 => (x"0e",x"4f",x"26",x"4b"),
   188 => (x"5d",x"5c",x"5b",x"5e"),
   189 => (x"ff",x"4d",x"71",x"0e"),
   190 => (x"49",x"75",x"4c",x"d4"),
   191 => (x"71",x"99",x"ff",x"c3"),
   192 => (x"c4",x"fe",x"c3",x"7c"),
   193 => (x"87",x"c8",x"05",x"bf"),
   194 => (x"c9",x"48",x"66",x"d0"),
   195 => (x"58",x"a6",x"d4",x"30"),
   196 => (x"d8",x"49",x"66",x"d0"),
   197 => (x"99",x"ff",x"c3",x"29"),
   198 => (x"66",x"d0",x"7c",x"71"),
   199 => (x"c3",x"29",x"d0",x"49"),
   200 => (x"7c",x"71",x"99",x"ff"),
   201 => (x"c8",x"49",x"66",x"d0"),
   202 => (x"99",x"ff",x"c3",x"29"),
   203 => (x"66",x"d0",x"7c",x"71"),
   204 => (x"99",x"ff",x"c3",x"49"),
   205 => (x"49",x"75",x"7c",x"71"),
   206 => (x"ff",x"c3",x"29",x"d0"),
   207 => (x"6c",x"7c",x"71",x"99"),
   208 => (x"ff",x"f0",x"c9",x"4b"),
   209 => (x"ab",x"ff",x"c3",x"4a"),
   210 => (x"49",x"87",x"cf",x"05"),
   211 => (x"4b",x"6c",x"7c",x"71"),
   212 => (x"c5",x"02",x"8a",x"c1"),
   213 => (x"02",x"ab",x"71",x"87"),
   214 => (x"48",x"73",x"87",x"f2"),
   215 => (x"4c",x"26",x"4d",x"26"),
   216 => (x"4f",x"26",x"4b",x"26"),
   217 => (x"ff",x"49",x"c0",x"1e"),
   218 => (x"ff",x"c3",x"48",x"d4"),
   219 => (x"c3",x"81",x"c1",x"78"),
   220 => (x"04",x"a9",x"b7",x"c8"),
   221 => (x"4f",x"26",x"87",x"f1"),
   222 => (x"5c",x"5b",x"5e",x"0e"),
   223 => (x"ff",x"c0",x"0e",x"5d"),
   224 => (x"4d",x"f7",x"c1",x"f0"),
   225 => (x"c0",x"c0",x"c0",x"c1"),
   226 => (x"ff",x"4b",x"c0",x"c0"),
   227 => (x"f8",x"c4",x"87",x"d6"),
   228 => (x"1e",x"c0",x"4c",x"df"),
   229 => (x"d6",x"fd",x"49",x"75"),
   230 => (x"c1",x"86",x"c4",x"87"),
   231 => (x"e5",x"c0",x"05",x"a8"),
   232 => (x"48",x"d4",x"ff",x"87"),
   233 => (x"73",x"78",x"ff",x"c3"),
   234 => (x"f0",x"e1",x"c0",x"1e"),
   235 => (x"fc",x"49",x"e9",x"c1"),
   236 => (x"86",x"c4",x"87",x"fd"),
   237 => (x"ca",x"05",x"98",x"70"),
   238 => (x"48",x"d4",x"ff",x"87"),
   239 => (x"c1",x"78",x"ff",x"c3"),
   240 => (x"fe",x"87",x"cb",x"48"),
   241 => (x"8c",x"c1",x"87",x"de"),
   242 => (x"87",x"c6",x"ff",x"05"),
   243 => (x"4d",x"26",x"48",x"c0"),
   244 => (x"4b",x"26",x"4c",x"26"),
   245 => (x"5e",x"0e",x"4f",x"26"),
   246 => (x"c0",x"0e",x"5c",x"5b"),
   247 => (x"c1",x"c1",x"f0",x"ff"),
   248 => (x"48",x"d4",x"ff",x"4c"),
   249 => (x"d3",x"78",x"ff",x"c3"),
   250 => (x"74",x"1e",x"c0",x"4b"),
   251 => (x"87",x"ff",x"fb",x"49"),
   252 => (x"98",x"70",x"86",x"c4"),
   253 => (x"ff",x"87",x"ca",x"05"),
   254 => (x"ff",x"c3",x"48",x"d4"),
   255 => (x"ca",x"48",x"c1",x"78"),
   256 => (x"87",x"e0",x"fd",x"87"),
   257 => (x"e0",x"05",x"8b",x"c1"),
   258 => (x"26",x"48",x"c0",x"87"),
   259 => (x"26",x"4b",x"26",x"4c"),
   260 => (x"5b",x"5e",x"0e",x"4f"),
   261 => (x"c3",x"0e",x"5d",x"5c"),
   262 => (x"d4",x"ff",x"4d",x"ff"),
   263 => (x"87",x"c4",x"fd",x"4b"),
   264 => (x"c0",x"1e",x"ea",x"c6"),
   265 => (x"c8",x"c1",x"f0",x"e1"),
   266 => (x"87",x"c3",x"fb",x"49"),
   267 => (x"a8",x"c1",x"86",x"c4"),
   268 => (x"fe",x"87",x"c8",x"02"),
   269 => (x"48",x"c0",x"87",x"e0"),
   270 => (x"fa",x"87",x"e2",x"c1"),
   271 => (x"49",x"70",x"87",x"c5"),
   272 => (x"99",x"ff",x"ff",x"cf"),
   273 => (x"02",x"a9",x"ea",x"c6"),
   274 => (x"c9",x"fe",x"87",x"c8"),
   275 => (x"c1",x"48",x"c0",x"87"),
   276 => (x"7b",x"75",x"87",x"cb"),
   277 => (x"fc",x"4c",x"f1",x"c0"),
   278 => (x"98",x"70",x"87",x"de"),
   279 => (x"87",x"ec",x"c0",x"02"),
   280 => (x"ff",x"c0",x"1e",x"c0"),
   281 => (x"49",x"fa",x"c1",x"f0"),
   282 => (x"c4",x"87",x"c4",x"fa"),
   283 => (x"05",x"98",x"70",x"86"),
   284 => (x"7b",x"75",x"87",x"da"),
   285 => (x"7b",x"75",x"49",x"6b"),
   286 => (x"7b",x"75",x"7b",x"75"),
   287 => (x"c0",x"c1",x"7b",x"75"),
   288 => (x"87",x"c4",x"02",x"99"),
   289 => (x"87",x"d5",x"48",x"c1"),
   290 => (x"87",x"d1",x"48",x"c0"),
   291 => (x"c4",x"05",x"ac",x"c2"),
   292 => (x"c8",x"48",x"c0",x"87"),
   293 => (x"05",x"8c",x"c1",x"87"),
   294 => (x"c0",x"87",x"fc",x"fe"),
   295 => (x"26",x"4d",x"26",x"48"),
   296 => (x"26",x"4b",x"26",x"4c"),
   297 => (x"5b",x"5e",x"0e",x"4f"),
   298 => (x"ff",x"0e",x"5d",x"5c"),
   299 => (x"e5",x"c0",x"4d",x"d0"),
   300 => (x"4c",x"c0",x"c1",x"d0"),
   301 => (x"48",x"c4",x"fe",x"c3"),
   302 => (x"4b",x"c7",x"78",x"c1"),
   303 => (x"e3",x"fa",x"7d",x"c2"),
   304 => (x"c0",x"7d",x"c3",x"87"),
   305 => (x"f8",x"49",x"74",x"1e"),
   306 => (x"86",x"c4",x"87",x"e5"),
   307 => (x"c1",x"05",x"a8",x"c1"),
   308 => (x"ab",x"c2",x"4b",x"87"),
   309 => (x"c0",x"87",x"c5",x"05"),
   310 => (x"87",x"f6",x"c0",x"48"),
   311 => (x"ff",x"05",x"8b",x"c1"),
   312 => (x"ec",x"fc",x"87",x"da"),
   313 => (x"c8",x"fe",x"c3",x"87"),
   314 => (x"05",x"98",x"70",x"58"),
   315 => (x"1e",x"c1",x"87",x"cd"),
   316 => (x"c1",x"f0",x"ff",x"c0"),
   317 => (x"f6",x"f7",x"49",x"d0"),
   318 => (x"ff",x"86",x"c4",x"87"),
   319 => (x"ff",x"c3",x"48",x"d4"),
   320 => (x"87",x"c3",x"c3",x"78"),
   321 => (x"58",x"cc",x"fe",x"c3"),
   322 => (x"d4",x"ff",x"7d",x"c2"),
   323 => (x"78",x"ff",x"c3",x"48"),
   324 => (x"4d",x"26",x"48",x"c1"),
   325 => (x"4b",x"26",x"4c",x"26"),
   326 => (x"5e",x"0e",x"4f",x"26"),
   327 => (x"0e",x"5d",x"5c",x"5b"),
   328 => (x"4b",x"71",x"86",x"fc"),
   329 => (x"c0",x"4c",x"d4",x"ff"),
   330 => (x"cd",x"ee",x"c5",x"7e"),
   331 => (x"ff",x"c3",x"4a",x"df"),
   332 => (x"c3",x"49",x"6c",x"7c"),
   333 => (x"c0",x"05",x"a9",x"fe"),
   334 => (x"4d",x"74",x"87",x"f8"),
   335 => (x"cc",x"02",x"9b",x"73"),
   336 => (x"1e",x"66",x"d4",x"87"),
   337 => (x"d1",x"f5",x"49",x"73"),
   338 => (x"d4",x"86",x"c4",x"87"),
   339 => (x"48",x"d0",x"ff",x"87"),
   340 => (x"d4",x"78",x"d1",x"c4"),
   341 => (x"ff",x"c3",x"4a",x"66"),
   342 => (x"05",x"8a",x"c1",x"7d"),
   343 => (x"a6",x"d8",x"87",x"f8"),
   344 => (x"7c",x"ff",x"c3",x"5a"),
   345 => (x"05",x"9b",x"73",x"7c"),
   346 => (x"d0",x"ff",x"87",x"c5"),
   347 => (x"c1",x"78",x"d0",x"48"),
   348 => (x"8a",x"c1",x"7e",x"4a"),
   349 => (x"87",x"f6",x"fe",x"05"),
   350 => (x"8e",x"fc",x"48",x"6e"),
   351 => (x"4c",x"26",x"4d",x"26"),
   352 => (x"4f",x"26",x"4b",x"26"),
   353 => (x"71",x"1e",x"73",x"1e"),
   354 => (x"ff",x"4b",x"c0",x"4a"),
   355 => (x"ff",x"c3",x"48",x"d4"),
   356 => (x"48",x"d0",x"ff",x"78"),
   357 => (x"ff",x"78",x"c3",x"c4"),
   358 => (x"ff",x"c3",x"48",x"d4"),
   359 => (x"c0",x"1e",x"72",x"78"),
   360 => (x"d1",x"c1",x"f0",x"ff"),
   361 => (x"87",x"c7",x"f5",x"49"),
   362 => (x"98",x"70",x"86",x"c4"),
   363 => (x"c8",x"87",x"d2",x"05"),
   364 => (x"66",x"cc",x"1e",x"c0"),
   365 => (x"87",x"e2",x"fd",x"49"),
   366 => (x"4b",x"70",x"86",x"c4"),
   367 => (x"c2",x"48",x"d0",x"ff"),
   368 => (x"26",x"48",x"73",x"78"),
   369 => (x"0e",x"4f",x"26",x"4b"),
   370 => (x"5d",x"5c",x"5b",x"5e"),
   371 => (x"c0",x"1e",x"c0",x"0e"),
   372 => (x"c9",x"c1",x"f0",x"ff"),
   373 => (x"87",x"d7",x"f4",x"49"),
   374 => (x"fe",x"c3",x"1e",x"d2"),
   375 => (x"f9",x"fc",x"49",x"cc"),
   376 => (x"c0",x"86",x"c8",x"87"),
   377 => (x"d2",x"84",x"c1",x"4c"),
   378 => (x"f8",x"04",x"ac",x"b7"),
   379 => (x"cc",x"fe",x"c3",x"87"),
   380 => (x"c3",x"49",x"bf",x"97"),
   381 => (x"c0",x"c1",x"99",x"c0"),
   382 => (x"e7",x"c0",x"05",x"a9"),
   383 => (x"d3",x"fe",x"c3",x"87"),
   384 => (x"d0",x"49",x"bf",x"97"),
   385 => (x"d4",x"fe",x"c3",x"31"),
   386 => (x"c8",x"4a",x"bf",x"97"),
   387 => (x"c3",x"b1",x"72",x"32"),
   388 => (x"bf",x"97",x"d5",x"fe"),
   389 => (x"4c",x"71",x"b1",x"4a"),
   390 => (x"ff",x"ff",x"ff",x"cf"),
   391 => (x"ca",x"84",x"c1",x"9c"),
   392 => (x"87",x"e7",x"c1",x"34"),
   393 => (x"97",x"d5",x"fe",x"c3"),
   394 => (x"31",x"c1",x"49",x"bf"),
   395 => (x"fe",x"c3",x"99",x"c6"),
   396 => (x"4a",x"bf",x"97",x"d6"),
   397 => (x"72",x"2a",x"b7",x"c7"),
   398 => (x"d1",x"fe",x"c3",x"b1"),
   399 => (x"4d",x"4a",x"bf",x"97"),
   400 => (x"fe",x"c3",x"9d",x"cf"),
   401 => (x"4a",x"bf",x"97",x"d2"),
   402 => (x"32",x"ca",x"9a",x"c3"),
   403 => (x"97",x"d3",x"fe",x"c3"),
   404 => (x"33",x"c2",x"4b",x"bf"),
   405 => (x"fe",x"c3",x"b2",x"73"),
   406 => (x"4b",x"bf",x"97",x"d4"),
   407 => (x"c6",x"9b",x"c0",x"c3"),
   408 => (x"b2",x"73",x"2b",x"b7"),
   409 => (x"48",x"c1",x"81",x"c2"),
   410 => (x"49",x"70",x"30",x"71"),
   411 => (x"30",x"75",x"48",x"c1"),
   412 => (x"4c",x"72",x"4d",x"70"),
   413 => (x"94",x"71",x"84",x"c1"),
   414 => (x"ad",x"b7",x"c0",x"c8"),
   415 => (x"c1",x"87",x"cc",x"06"),
   416 => (x"c8",x"2d",x"b7",x"34"),
   417 => (x"01",x"ad",x"b7",x"c0"),
   418 => (x"74",x"87",x"f4",x"ff"),
   419 => (x"26",x"4d",x"26",x"48"),
   420 => (x"26",x"4b",x"26",x"4c"),
   421 => (x"5b",x"5e",x"0e",x"4f"),
   422 => (x"f8",x"0e",x"5d",x"5c"),
   423 => (x"f4",x"c6",x"c4",x"86"),
   424 => (x"c3",x"78",x"c0",x"48"),
   425 => (x"c0",x"1e",x"ec",x"fe"),
   426 => (x"87",x"d8",x"fb",x"49"),
   427 => (x"98",x"70",x"86",x"c4"),
   428 => (x"c0",x"87",x"c5",x"05"),
   429 => (x"87",x"ce",x"c9",x"48"),
   430 => (x"7e",x"c1",x"4d",x"c0"),
   431 => (x"bf",x"e0",x"fe",x"c0"),
   432 => (x"e2",x"ff",x"c3",x"49"),
   433 => (x"4b",x"c8",x"71",x"4a"),
   434 => (x"70",x"87",x"f0",x"e6"),
   435 => (x"87",x"c2",x"05",x"98"),
   436 => (x"fe",x"c0",x"7e",x"c0"),
   437 => (x"c3",x"49",x"bf",x"dc"),
   438 => (x"71",x"4a",x"fe",x"ff"),
   439 => (x"da",x"e6",x"4b",x"c8"),
   440 => (x"05",x"98",x"70",x"87"),
   441 => (x"7e",x"c0",x"87",x"c2"),
   442 => (x"fd",x"c0",x"02",x"6e"),
   443 => (x"f2",x"c5",x"c4",x"87"),
   444 => (x"c6",x"c4",x"4d",x"bf"),
   445 => (x"7e",x"bf",x"9f",x"ea"),
   446 => (x"ea",x"d6",x"c5",x"48"),
   447 => (x"87",x"c7",x"05",x"a8"),
   448 => (x"bf",x"f2",x"c5",x"c4"),
   449 => (x"6e",x"87",x"ce",x"4d"),
   450 => (x"d5",x"e9",x"ca",x"48"),
   451 => (x"87",x"c5",x"02",x"a8"),
   452 => (x"f1",x"c7",x"48",x"c0"),
   453 => (x"ec",x"fe",x"c3",x"87"),
   454 => (x"f9",x"49",x"75",x"1e"),
   455 => (x"86",x"c4",x"87",x"e6"),
   456 => (x"c5",x"05",x"98",x"70"),
   457 => (x"c7",x"48",x"c0",x"87"),
   458 => (x"fe",x"c0",x"87",x"dc"),
   459 => (x"c3",x"49",x"bf",x"dc"),
   460 => (x"71",x"4a",x"fe",x"ff"),
   461 => (x"c2",x"e5",x"4b",x"c8"),
   462 => (x"05",x"98",x"70",x"87"),
   463 => (x"c6",x"c4",x"87",x"c8"),
   464 => (x"78",x"c1",x"48",x"f4"),
   465 => (x"fe",x"c0",x"87",x"da"),
   466 => (x"c3",x"49",x"bf",x"e0"),
   467 => (x"71",x"4a",x"e2",x"ff"),
   468 => (x"e6",x"e4",x"4b",x"c8"),
   469 => (x"02",x"98",x"70",x"87"),
   470 => (x"c0",x"87",x"c5",x"c0"),
   471 => (x"87",x"e6",x"c6",x"48"),
   472 => (x"97",x"ea",x"c6",x"c4"),
   473 => (x"d5",x"c1",x"49",x"bf"),
   474 => (x"cd",x"c0",x"05",x"a9"),
   475 => (x"eb",x"c6",x"c4",x"87"),
   476 => (x"c2",x"49",x"bf",x"97"),
   477 => (x"c0",x"02",x"a9",x"ea"),
   478 => (x"48",x"c0",x"87",x"c5"),
   479 => (x"c3",x"87",x"c7",x"c6"),
   480 => (x"bf",x"97",x"ec",x"fe"),
   481 => (x"e9",x"c3",x"48",x"7e"),
   482 => (x"ce",x"c0",x"02",x"a8"),
   483 => (x"c3",x"48",x"6e",x"87"),
   484 => (x"c0",x"02",x"a8",x"eb"),
   485 => (x"48",x"c0",x"87",x"c5"),
   486 => (x"c3",x"87",x"eb",x"c5"),
   487 => (x"bf",x"97",x"f7",x"fe"),
   488 => (x"c0",x"05",x"99",x"49"),
   489 => (x"fe",x"c3",x"87",x"cc"),
   490 => (x"49",x"bf",x"97",x"f8"),
   491 => (x"c0",x"02",x"a9",x"c2"),
   492 => (x"48",x"c0",x"87",x"c5"),
   493 => (x"c3",x"87",x"cf",x"c5"),
   494 => (x"bf",x"97",x"f9",x"fe"),
   495 => (x"f0",x"c6",x"c4",x"48"),
   496 => (x"48",x"4c",x"70",x"58"),
   497 => (x"c6",x"c4",x"88",x"c1"),
   498 => (x"fe",x"c3",x"58",x"f4"),
   499 => (x"49",x"bf",x"97",x"fa"),
   500 => (x"fe",x"c3",x"81",x"75"),
   501 => (x"4a",x"bf",x"97",x"fb"),
   502 => (x"a1",x"72",x"32",x"c8"),
   503 => (x"c4",x"cb",x"c4",x"7e"),
   504 => (x"c3",x"78",x"6e",x"48"),
   505 => (x"bf",x"97",x"fc",x"fe"),
   506 => (x"58",x"a6",x"c8",x"48"),
   507 => (x"bf",x"f4",x"c6",x"c4"),
   508 => (x"87",x"d4",x"c2",x"02"),
   509 => (x"bf",x"dc",x"fe",x"c0"),
   510 => (x"fe",x"ff",x"c3",x"49"),
   511 => (x"4b",x"c8",x"71",x"4a"),
   512 => (x"70",x"87",x"f8",x"e1"),
   513 => (x"c5",x"c0",x"02",x"98"),
   514 => (x"c3",x"48",x"c0",x"87"),
   515 => (x"c6",x"c4",x"87",x"f8"),
   516 => (x"c4",x"4c",x"bf",x"ec"),
   517 => (x"c3",x"5c",x"d8",x"cb"),
   518 => (x"bf",x"97",x"d1",x"ff"),
   519 => (x"c3",x"31",x"c8",x"49"),
   520 => (x"bf",x"97",x"d0",x"ff"),
   521 => (x"c3",x"49",x"a1",x"4a"),
   522 => (x"bf",x"97",x"d2",x"ff"),
   523 => (x"72",x"32",x"d0",x"4a"),
   524 => (x"ff",x"c3",x"49",x"a1"),
   525 => (x"4a",x"bf",x"97",x"d3"),
   526 => (x"a1",x"72",x"32",x"d8"),
   527 => (x"91",x"66",x"c4",x"49"),
   528 => (x"bf",x"c4",x"cb",x"c4"),
   529 => (x"cc",x"cb",x"c4",x"81"),
   530 => (x"d9",x"ff",x"c3",x"59"),
   531 => (x"c8",x"4a",x"bf",x"97"),
   532 => (x"d8",x"ff",x"c3",x"32"),
   533 => (x"a2",x"4b",x"bf",x"97"),
   534 => (x"da",x"ff",x"c3",x"4a"),
   535 => (x"d0",x"4b",x"bf",x"97"),
   536 => (x"4a",x"a2",x"73",x"33"),
   537 => (x"97",x"db",x"ff",x"c3"),
   538 => (x"9b",x"cf",x"4b",x"bf"),
   539 => (x"a2",x"73",x"33",x"d8"),
   540 => (x"d0",x"cb",x"c4",x"4a"),
   541 => (x"cc",x"cb",x"c4",x"5a"),
   542 => (x"8a",x"c2",x"4a",x"bf"),
   543 => (x"cb",x"c4",x"92",x"74"),
   544 => (x"a1",x"72",x"48",x"d0"),
   545 => (x"87",x"ca",x"c1",x"78"),
   546 => (x"97",x"fe",x"fe",x"c3"),
   547 => (x"31",x"c8",x"49",x"bf"),
   548 => (x"97",x"fd",x"fe",x"c3"),
   549 => (x"49",x"a1",x"4a",x"bf"),
   550 => (x"59",x"fc",x"c6",x"c4"),
   551 => (x"bf",x"f8",x"c6",x"c4"),
   552 => (x"c7",x"31",x"c5",x"49"),
   553 => (x"29",x"c9",x"81",x"ff"),
   554 => (x"59",x"d8",x"cb",x"c4"),
   555 => (x"97",x"c3",x"ff",x"c3"),
   556 => (x"32",x"c8",x"4a",x"bf"),
   557 => (x"97",x"c2",x"ff",x"c3"),
   558 => (x"4a",x"a2",x"4b",x"bf"),
   559 => (x"6e",x"92",x"66",x"c4"),
   560 => (x"d4",x"cb",x"c4",x"82"),
   561 => (x"cc",x"cb",x"c4",x"5a"),
   562 => (x"c4",x"78",x"c0",x"48"),
   563 => (x"72",x"48",x"c8",x"cb"),
   564 => (x"cb",x"c4",x"78",x"a1"),
   565 => (x"cb",x"c4",x"48",x"d8"),
   566 => (x"c4",x"78",x"bf",x"cc"),
   567 => (x"c4",x"48",x"dc",x"cb"),
   568 => (x"78",x"bf",x"d0",x"cb"),
   569 => (x"bf",x"f4",x"c6",x"c4"),
   570 => (x"87",x"c9",x"c0",x"02"),
   571 => (x"30",x"c4",x"48",x"74"),
   572 => (x"c9",x"c0",x"7e",x"70"),
   573 => (x"d4",x"cb",x"c4",x"87"),
   574 => (x"30",x"c4",x"48",x"bf"),
   575 => (x"c6",x"c4",x"7e",x"70"),
   576 => (x"78",x"6e",x"48",x"f8"),
   577 => (x"8e",x"f8",x"48",x"c1"),
   578 => (x"4c",x"26",x"4d",x"26"),
   579 => (x"4f",x"26",x"4b",x"26"),
   580 => (x"5c",x"5b",x"5e",x"0e"),
   581 => (x"4a",x"71",x"0e",x"5d"),
   582 => (x"bf",x"f4",x"c6",x"c4"),
   583 => (x"72",x"87",x"cb",x"02"),
   584 => (x"72",x"2b",x"c7",x"4b"),
   585 => (x"9c",x"ff",x"c1",x"4c"),
   586 => (x"4b",x"72",x"87",x"c9"),
   587 => (x"4c",x"72",x"2b",x"c8"),
   588 => (x"c4",x"9c",x"ff",x"c3"),
   589 => (x"83",x"bf",x"c4",x"cb"),
   590 => (x"bf",x"d8",x"fe",x"c0"),
   591 => (x"87",x"d9",x"02",x"ab"),
   592 => (x"5b",x"dc",x"fe",x"c0"),
   593 => (x"1e",x"ec",x"fe",x"c3"),
   594 => (x"f7",x"f0",x"49",x"73"),
   595 => (x"70",x"86",x"c4",x"87"),
   596 => (x"87",x"c5",x"05",x"98"),
   597 => (x"e6",x"c0",x"48",x"c0"),
   598 => (x"f4",x"c6",x"c4",x"87"),
   599 => (x"87",x"d2",x"02",x"bf"),
   600 => (x"91",x"c4",x"49",x"74"),
   601 => (x"81",x"ec",x"fe",x"c3"),
   602 => (x"ff",x"cf",x"4d",x"69"),
   603 => (x"9d",x"ff",x"ff",x"ff"),
   604 => (x"49",x"74",x"87",x"cb"),
   605 => (x"fe",x"c3",x"91",x"c2"),
   606 => (x"69",x"9f",x"81",x"ec"),
   607 => (x"26",x"48",x"75",x"4d"),
   608 => (x"26",x"4c",x"26",x"4d"),
   609 => (x"0e",x"4f",x"26",x"4b"),
   610 => (x"5d",x"5c",x"5b",x"5e"),
   611 => (x"cc",x"86",x"f4",x"0e"),
   612 => (x"66",x"c8",x"59",x"a6"),
   613 => (x"c0",x"87",x"c5",x"05"),
   614 => (x"87",x"c8",x"c3",x"48"),
   615 => (x"c8",x"48",x"66",x"c8"),
   616 => (x"6e",x"7e",x"70",x"80"),
   617 => (x"dc",x"78",x"c0",x"48"),
   618 => (x"87",x"c7",x"02",x"66"),
   619 => (x"bf",x"97",x"66",x"dc"),
   620 => (x"c0",x"87",x"c5",x"05"),
   621 => (x"87",x"ec",x"c2",x"48"),
   622 => (x"49",x"c1",x"1e",x"c0"),
   623 => (x"c4",x"87",x"db",x"cf"),
   624 => (x"9c",x"4c",x"70",x"86"),
   625 => (x"87",x"fc",x"c0",x"02"),
   626 => (x"4a",x"fc",x"c6",x"c4"),
   627 => (x"ff",x"49",x"66",x"dc"),
   628 => (x"70",x"87",x"cd",x"da"),
   629 => (x"eb",x"c0",x"02",x"98"),
   630 => (x"dc",x"4a",x"74",x"87"),
   631 => (x"4b",x"cb",x"49",x"66"),
   632 => (x"87",x"f1",x"da",x"ff"),
   633 => (x"db",x"02",x"98",x"70"),
   634 => (x"74",x"1e",x"c0",x"87"),
   635 => (x"87",x"c4",x"02",x"9c"),
   636 => (x"87",x"c2",x"4d",x"c0"),
   637 => (x"49",x"75",x"4d",x"c1"),
   638 => (x"c4",x"87",x"df",x"ce"),
   639 => (x"9c",x"4c",x"70",x"86"),
   640 => (x"87",x"c4",x"ff",x"05"),
   641 => (x"c1",x"02",x"9c",x"74"),
   642 => (x"a4",x"dc",x"87",x"d8"),
   643 => (x"69",x"48",x"6e",x"49"),
   644 => (x"49",x"a4",x"da",x"78"),
   645 => (x"c4",x"48",x"66",x"c8"),
   646 => (x"58",x"a6",x"c8",x"80"),
   647 => (x"c4",x"48",x"69",x"9f"),
   648 => (x"c4",x"78",x"08",x"66"),
   649 => (x"02",x"bf",x"f4",x"c6"),
   650 => (x"a4",x"d4",x"87",x"d2"),
   651 => (x"49",x"69",x"9f",x"49"),
   652 => (x"99",x"ff",x"ff",x"c0"),
   653 => (x"30",x"d0",x"48",x"71"),
   654 => (x"87",x"c2",x"7e",x"70"),
   655 => (x"49",x"6e",x"7e",x"c0"),
   656 => (x"bf",x"66",x"c4",x"48"),
   657 => (x"08",x"66",x"c4",x"80"),
   658 => (x"48",x"66",x"c8",x"78"),
   659 => (x"66",x"c8",x"78",x"c0"),
   660 => (x"c4",x"81",x"cc",x"49"),
   661 => (x"c8",x"79",x"bf",x"66"),
   662 => (x"81",x"d0",x"49",x"66"),
   663 => (x"48",x"c1",x"79",x"c0"),
   664 => (x"48",x"c0",x"87",x"c2"),
   665 => (x"4d",x"26",x"8e",x"f4"),
   666 => (x"4b",x"26",x"4c",x"26"),
   667 => (x"5e",x"0e",x"4f",x"26"),
   668 => (x"0e",x"5d",x"5c",x"5b"),
   669 => (x"02",x"9c",x"4c",x"71"),
   670 => (x"c8",x"87",x"ca",x"c1"),
   671 => (x"02",x"69",x"49",x"a4"),
   672 => (x"d0",x"87",x"c2",x"c1"),
   673 => (x"49",x"6c",x"4a",x"66"),
   674 => (x"5a",x"a6",x"d4",x"82"),
   675 => (x"b9",x"4d",x"66",x"d0"),
   676 => (x"bf",x"f0",x"c6",x"c4"),
   677 => (x"72",x"ba",x"ff",x"4a"),
   678 => (x"02",x"99",x"71",x"99"),
   679 => (x"c4",x"87",x"e4",x"c0"),
   680 => (x"49",x"6b",x"4b",x"a4"),
   681 => (x"70",x"87",x"e9",x"f9"),
   682 => (x"ec",x"c6",x"c4",x"7b"),
   683 => (x"81",x"6c",x"49",x"bf"),
   684 => (x"b9",x"75",x"7c",x"71"),
   685 => (x"bf",x"f0",x"c6",x"c4"),
   686 => (x"72",x"ba",x"ff",x"4a"),
   687 => (x"05",x"99",x"71",x"99"),
   688 => (x"75",x"87",x"dc",x"ff"),
   689 => (x"26",x"4d",x"26",x"7c"),
   690 => (x"26",x"4b",x"26",x"4c"),
   691 => (x"1e",x"73",x"1e",x"4f"),
   692 => (x"02",x"9b",x"4b",x"71"),
   693 => (x"a3",x"c8",x"87",x"c7"),
   694 => (x"c5",x"05",x"69",x"49"),
   695 => (x"c0",x"48",x"c0",x"87"),
   696 => (x"cb",x"c4",x"87",x"f7"),
   697 => (x"c4",x"4a",x"bf",x"c8"),
   698 => (x"49",x"69",x"49",x"a3"),
   699 => (x"c6",x"c4",x"89",x"c2"),
   700 => (x"71",x"91",x"bf",x"ec"),
   701 => (x"c6",x"c4",x"4a",x"a2"),
   702 => (x"6b",x"49",x"bf",x"f0"),
   703 => (x"4a",x"a2",x"71",x"99"),
   704 => (x"5a",x"dc",x"fe",x"c0"),
   705 => (x"72",x"1e",x"66",x"c8"),
   706 => (x"87",x"f8",x"e9",x"49"),
   707 => (x"98",x"70",x"86",x"c4"),
   708 => (x"c0",x"87",x"c4",x"05"),
   709 => (x"c1",x"87",x"c2",x"48"),
   710 => (x"26",x"4b",x"26",x"48"),
   711 => (x"5b",x"5e",x"0e",x"4f"),
   712 => (x"fc",x"0e",x"5d",x"5c"),
   713 => (x"d4",x"4b",x"71",x"86"),
   714 => (x"9b",x"73",x"4d",x"66"),
   715 => (x"87",x"cc",x"c1",x"02"),
   716 => (x"69",x"49",x"a3",x"c8"),
   717 => (x"87",x"c4",x"c1",x"02"),
   718 => (x"c4",x"4c",x"a3",x"d0"),
   719 => (x"49",x"bf",x"f0",x"c6"),
   720 => (x"4a",x"6c",x"b9",x"ff"),
   721 => (x"66",x"d4",x"7e",x"99"),
   722 => (x"87",x"cd",x"06",x"a9"),
   723 => (x"cc",x"7c",x"7b",x"c0"),
   724 => (x"a3",x"c4",x"4a",x"a3"),
   725 => (x"ca",x"79",x"6a",x"49"),
   726 => (x"f8",x"49",x"72",x"87"),
   727 => (x"66",x"d4",x"99",x"c0"),
   728 => (x"75",x"8d",x"71",x"4d"),
   729 => (x"71",x"29",x"c9",x"49"),
   730 => (x"fc",x"49",x"73",x"1e"),
   731 => (x"fe",x"c3",x"87",x"c0"),
   732 => (x"49",x"73",x"1e",x"ec"),
   733 => (x"c8",x"87",x"d6",x"fd"),
   734 => (x"7c",x"66",x"d4",x"86"),
   735 => (x"4d",x"26",x"8e",x"fc"),
   736 => (x"4b",x"26",x"4c",x"26"),
   737 => (x"5e",x"0e",x"4f",x"26"),
   738 => (x"0e",x"5d",x"5c",x"5b"),
   739 => (x"a6",x"d0",x"86",x"f0"),
   740 => (x"66",x"e0",x"c0",x"59"),
   741 => (x"66",x"e4",x"c0",x"4c"),
   742 => (x"02",x"66",x"cc",x"4b"),
   743 => (x"c8",x"48",x"87",x"ca"),
   744 => (x"6e",x"7e",x"70",x"80"),
   745 => (x"87",x"c5",x"05",x"bf"),
   746 => (x"ec",x"c3",x"48",x"c0"),
   747 => (x"4d",x"66",x"cc",x"87"),
   748 => (x"49",x"73",x"85",x"d0"),
   749 => (x"6d",x"48",x"a6",x"c4"),
   750 => (x"81",x"66",x"c4",x"78"),
   751 => (x"bf",x"6e",x"80",x"c4"),
   752 => (x"a9",x"66",x"c8",x"78"),
   753 => (x"49",x"87",x"c6",x"06"),
   754 => (x"71",x"89",x"66",x"c4"),
   755 => (x"ab",x"b7",x"c0",x"4b"),
   756 => (x"48",x"87",x"c4",x"01"),
   757 => (x"c4",x"87",x"c2",x"c3"),
   758 => (x"ff",x"c7",x"48",x"66"),
   759 => (x"6e",x"7e",x"70",x"98"),
   760 => (x"87",x"cd",x"c1",x"02"),
   761 => (x"6e",x"49",x"c0",x"c8"),
   762 => (x"59",x"a6",x"cc",x"89"),
   763 => (x"4a",x"ec",x"fe",x"c3"),
   764 => (x"66",x"c8",x"82",x"6e"),
   765 => (x"c3",x"03",x"ab",x"b7"),
   766 => (x"5b",x"a6",x"cc",x"87"),
   767 => (x"48",x"49",x"66",x"c8"),
   768 => (x"70",x"80",x"66",x"c4"),
   769 => (x"8b",x"66",x"c8",x"7d"),
   770 => (x"88",x"c1",x"48",x"49"),
   771 => (x"71",x"58",x"a6",x"cc"),
   772 => (x"87",x"d3",x"02",x"99"),
   773 => (x"c1",x"7c",x"97",x"12"),
   774 => (x"49",x"66",x"c8",x"84"),
   775 => (x"cc",x"88",x"c1",x"48"),
   776 => (x"99",x"71",x"58",x"a6"),
   777 => (x"c1",x"87",x"ed",x"05"),
   778 => (x"49",x"66",x"d0",x"1e"),
   779 => (x"c4",x"87",x"ff",x"f8"),
   780 => (x"ab",x"b7",x"c0",x"86"),
   781 => (x"87",x"df",x"c1",x"06"),
   782 => (x"ab",x"b7",x"ff",x"c7"),
   783 => (x"87",x"e2",x"c0",x"06"),
   784 => (x"66",x"d0",x"1e",x"74"),
   785 => (x"87",x"c5",x"fa",x"49"),
   786 => (x"6d",x"84",x"c0",x"c8"),
   787 => (x"80",x"c0",x"c8",x"48"),
   788 => (x"c0",x"c8",x"7d",x"70"),
   789 => (x"d4",x"1e",x"c1",x"8b"),
   790 => (x"d1",x"f8",x"49",x"66"),
   791 => (x"c0",x"86",x"c8",x"87"),
   792 => (x"fe",x"c3",x"87",x"ee"),
   793 => (x"66",x"d0",x"1e",x"ec"),
   794 => (x"87",x"e1",x"f9",x"49"),
   795 => (x"fe",x"c3",x"86",x"c4"),
   796 => (x"49",x"73",x"4a",x"ec"),
   797 => (x"70",x"80",x"6d",x"48"),
   798 => (x"c1",x"49",x"73",x"7d"),
   799 => (x"02",x"99",x"71",x"8b"),
   800 => (x"97",x"12",x"87",x"ce"),
   801 => (x"73",x"84",x"c1",x"7c"),
   802 => (x"71",x"8b",x"c1",x"49"),
   803 => (x"87",x"f2",x"05",x"99"),
   804 => (x"01",x"ab",x"b7",x"c0"),
   805 => (x"c1",x"87",x"e1",x"fe"),
   806 => (x"26",x"8e",x"f0",x"48"),
   807 => (x"26",x"4c",x"26",x"4d"),
   808 => (x"0e",x"4f",x"26",x"4b"),
   809 => (x"5d",x"5c",x"5b",x"5e"),
   810 => (x"9b",x"4b",x"71",x"0e"),
   811 => (x"c8",x"87",x"c7",x"02"),
   812 => (x"05",x"6d",x"4d",x"a3"),
   813 => (x"48",x"ff",x"87",x"c5"),
   814 => (x"d0",x"87",x"fd",x"c0"),
   815 => (x"49",x"6c",x"4c",x"a3"),
   816 => (x"05",x"99",x"ff",x"c7"),
   817 => (x"02",x"6c",x"87",x"d8"),
   818 => (x"1e",x"c1",x"87",x"c9"),
   819 => (x"dd",x"f6",x"49",x"73"),
   820 => (x"c3",x"86",x"c4",x"87"),
   821 => (x"73",x"1e",x"ec",x"fe"),
   822 => (x"87",x"f1",x"f7",x"49"),
   823 => (x"4a",x"6c",x"86",x"c4"),
   824 => (x"c4",x"04",x"aa",x"6d"),
   825 => (x"cf",x"48",x"ff",x"87"),
   826 => (x"7c",x"a2",x"c1",x"87"),
   827 => (x"ff",x"c7",x"49",x"72"),
   828 => (x"ec",x"fe",x"c3",x"99"),
   829 => (x"48",x"69",x"97",x"81"),
   830 => (x"4c",x"26",x"4d",x"26"),
   831 => (x"4f",x"26",x"4b",x"26"),
   832 => (x"71",x"1e",x"73",x"1e"),
   833 => (x"c0",x"02",x"9b",x"4b"),
   834 => (x"cb",x"c4",x"87",x"e4"),
   835 => (x"4a",x"73",x"5b",x"dc"),
   836 => (x"c6",x"c4",x"8a",x"c2"),
   837 => (x"92",x"49",x"bf",x"ec"),
   838 => (x"bf",x"c8",x"cb",x"c4"),
   839 => (x"c4",x"80",x"72",x"48"),
   840 => (x"71",x"58",x"e0",x"cb"),
   841 => (x"c4",x"30",x"c4",x"48"),
   842 => (x"c0",x"58",x"fc",x"c6"),
   843 => (x"cb",x"c4",x"87",x"ed"),
   844 => (x"cb",x"c4",x"48",x"d8"),
   845 => (x"c4",x"78",x"bf",x"cc"),
   846 => (x"c4",x"48",x"dc",x"cb"),
   847 => (x"78",x"bf",x"d0",x"cb"),
   848 => (x"bf",x"f4",x"c6",x"c4"),
   849 => (x"c4",x"87",x"c9",x"02"),
   850 => (x"49",x"bf",x"ec",x"c6"),
   851 => (x"87",x"c7",x"31",x"c4"),
   852 => (x"bf",x"d4",x"cb",x"c4"),
   853 => (x"c4",x"31",x"c4",x"49"),
   854 => (x"26",x"59",x"fc",x"c6"),
   855 => (x"0e",x"4f",x"26",x"4b"),
   856 => (x"0e",x"5c",x"5b",x"5e"),
   857 => (x"4b",x"c0",x"4a",x"71"),
   858 => (x"c0",x"02",x"9a",x"72"),
   859 => (x"a2",x"da",x"87",x"e1"),
   860 => (x"4b",x"69",x"9f",x"49"),
   861 => (x"bf",x"f4",x"c6",x"c4"),
   862 => (x"d4",x"87",x"cf",x"02"),
   863 => (x"69",x"9f",x"49",x"a2"),
   864 => (x"ff",x"c0",x"4c",x"49"),
   865 => (x"34",x"d0",x"9c",x"ff"),
   866 => (x"4c",x"c0",x"87",x"c2"),
   867 => (x"73",x"b3",x"49",x"74"),
   868 => (x"87",x"ec",x"fd",x"49"),
   869 => (x"4b",x"26",x"4c",x"26"),
   870 => (x"5e",x"0e",x"4f",x"26"),
   871 => (x"0e",x"5d",x"5c",x"5b"),
   872 => (x"a6",x"c8",x"86",x"f0"),
   873 => (x"ff",x"ff",x"cf",x"59"),
   874 => (x"c0",x"4c",x"f8",x"ff"),
   875 => (x"02",x"66",x"c4",x"7e"),
   876 => (x"fe",x"c3",x"87",x"d8"),
   877 => (x"78",x"c0",x"48",x"e8"),
   878 => (x"48",x"e0",x"fe",x"c3"),
   879 => (x"bf",x"dc",x"cb",x"c4"),
   880 => (x"e4",x"fe",x"c3",x"78"),
   881 => (x"d8",x"cb",x"c4",x"48"),
   882 => (x"c7",x"c4",x"78",x"bf"),
   883 => (x"50",x"c0",x"48",x"c9"),
   884 => (x"bf",x"f8",x"c6",x"c4"),
   885 => (x"e8",x"fe",x"c3",x"49"),
   886 => (x"aa",x"71",x"4a",x"bf"),
   887 => (x"87",x"cc",x"c4",x"03"),
   888 => (x"99",x"cf",x"49",x"72"),
   889 => (x"87",x"ea",x"c0",x"05"),
   890 => (x"48",x"d8",x"fe",x"c0"),
   891 => (x"bf",x"e0",x"fe",x"c3"),
   892 => (x"ec",x"fe",x"c3",x"78"),
   893 => (x"e0",x"fe",x"c3",x"1e"),
   894 => (x"fe",x"c3",x"49",x"bf"),
   895 => (x"a1",x"c1",x"48",x"e0"),
   896 => (x"dd",x"ff",x"71",x"78"),
   897 => (x"86",x"c4",x"87",x"fe"),
   898 => (x"48",x"d4",x"fe",x"c0"),
   899 => (x"78",x"ec",x"fe",x"c3"),
   900 => (x"fe",x"c0",x"87",x"cc"),
   901 => (x"c0",x"48",x"bf",x"d4"),
   902 => (x"fe",x"c0",x"80",x"e0"),
   903 => (x"fe",x"c3",x"58",x"d8"),
   904 => (x"c1",x"48",x"bf",x"e8"),
   905 => (x"ec",x"fe",x"c3",x"80"),
   906 => (x"0f",x"94",x"27",x"58"),
   907 => (x"97",x"bf",x"00",x"00"),
   908 => (x"02",x"9d",x"4d",x"bf"),
   909 => (x"c3",x"87",x"e5",x"c2"),
   910 => (x"c2",x"02",x"ad",x"e5"),
   911 => (x"fe",x"c0",x"87",x"de"),
   912 => (x"cb",x"4b",x"bf",x"d4"),
   913 => (x"4c",x"11",x"49",x"a3"),
   914 => (x"c1",x"05",x"ac",x"cf"),
   915 => (x"49",x"75",x"87",x"d2"),
   916 => (x"89",x"c1",x"99",x"df"),
   917 => (x"c6",x"c4",x"91",x"cd"),
   918 => (x"a3",x"c1",x"81",x"fc"),
   919 => (x"c3",x"51",x"12",x"4a"),
   920 => (x"51",x"12",x"4a",x"a3"),
   921 => (x"12",x"4a",x"a3",x"c5"),
   922 => (x"4a",x"a3",x"c7",x"51"),
   923 => (x"a3",x"c9",x"51",x"12"),
   924 => (x"ce",x"51",x"12",x"4a"),
   925 => (x"51",x"12",x"4a",x"a3"),
   926 => (x"12",x"4a",x"a3",x"d0"),
   927 => (x"4a",x"a3",x"d2",x"51"),
   928 => (x"a3",x"d4",x"51",x"12"),
   929 => (x"d6",x"51",x"12",x"4a"),
   930 => (x"51",x"12",x"4a",x"a3"),
   931 => (x"12",x"4a",x"a3",x"d8"),
   932 => (x"4a",x"a3",x"dc",x"51"),
   933 => (x"a3",x"de",x"51",x"12"),
   934 => (x"c1",x"51",x"12",x"4a"),
   935 => (x"87",x"fc",x"c0",x"7e"),
   936 => (x"99",x"c8",x"49",x"74"),
   937 => (x"87",x"ed",x"c0",x"05"),
   938 => (x"99",x"d0",x"49",x"74"),
   939 => (x"c0",x"87",x"d3",x"05"),
   940 => (x"c0",x"02",x"66",x"e0"),
   941 => (x"49",x"73",x"87",x"cc"),
   942 => (x"0f",x"66",x"e0",x"c0"),
   943 => (x"c0",x"02",x"98",x"70"),
   944 => (x"05",x"6e",x"87",x"d3"),
   945 => (x"c4",x"87",x"c6",x"c0"),
   946 => (x"c0",x"48",x"fc",x"c6"),
   947 => (x"d4",x"fe",x"c0",x"50"),
   948 => (x"ed",x"c2",x"48",x"bf"),
   949 => (x"c9",x"c7",x"c4",x"87"),
   950 => (x"7e",x"50",x"c0",x"48"),
   951 => (x"bf",x"f8",x"c6",x"c4"),
   952 => (x"e8",x"fe",x"c3",x"49"),
   953 => (x"aa",x"71",x"4a",x"bf"),
   954 => (x"87",x"f4",x"fb",x"04"),
   955 => (x"ff",x"ff",x"ff",x"cf"),
   956 => (x"cb",x"c4",x"4c",x"f8"),
   957 => (x"c0",x"05",x"bf",x"dc"),
   958 => (x"c6",x"c4",x"87",x"c8"),
   959 => (x"c1",x"02",x"bf",x"f4"),
   960 => (x"fe",x"c3",x"87",x"fe"),
   961 => (x"e8",x"49",x"bf",x"e4"),
   962 => (x"49",x"70",x"87",x"c6"),
   963 => (x"59",x"e8",x"fe",x"c3"),
   964 => (x"c3",x"48",x"a6",x"c4"),
   965 => (x"78",x"bf",x"e4",x"fe"),
   966 => (x"bf",x"f4",x"c6",x"c4"),
   967 => (x"87",x"db",x"c0",x"02"),
   968 => (x"74",x"49",x"66",x"c4"),
   969 => (x"02",x"a9",x"74",x"99"),
   970 => (x"c8",x"87",x"c8",x"c0"),
   971 => (x"78",x"c0",x"48",x"a6"),
   972 => (x"c8",x"87",x"e7",x"c0"),
   973 => (x"78",x"c1",x"48",x"a6"),
   974 => (x"c4",x"87",x"df",x"c0"),
   975 => (x"ff",x"cf",x"49",x"66"),
   976 => (x"02",x"a9",x"99",x"f8"),
   977 => (x"cc",x"87",x"c8",x"c0"),
   978 => (x"78",x"c0",x"48",x"a6"),
   979 => (x"cc",x"87",x"c5",x"c0"),
   980 => (x"78",x"c1",x"48",x"a6"),
   981 => (x"cc",x"48",x"a6",x"c8"),
   982 => (x"66",x"c8",x"78",x"66"),
   983 => (x"87",x"e0",x"c0",x"05"),
   984 => (x"c2",x"49",x"66",x"c4"),
   985 => (x"ec",x"c6",x"c4",x"89"),
   986 => (x"c4",x"91",x"4a",x"bf"),
   987 => (x"4a",x"bf",x"c8",x"cb"),
   988 => (x"48",x"e0",x"fe",x"c3"),
   989 => (x"c3",x"78",x"a1",x"72"),
   990 => (x"c0",x"48",x"e8",x"fe"),
   991 => (x"87",x"d0",x"f9",x"78"),
   992 => (x"ff",x"cf",x"48",x"c0"),
   993 => (x"4c",x"f8",x"ff",x"ff"),
   994 => (x"4d",x"26",x"8e",x"f0"),
   995 => (x"4b",x"26",x"4c",x"26"),
   996 => (x"00",x"00",x"4f",x"26"),
   997 => (x"00",x"00",x"00",x"00"),
   998 => (x"ff",x"ff",x"ff",x"ff"),
   999 => (x"00",x"00",x"0f",x"a4"),
  1000 => (x"00",x"00",x"0f",x"b0"),
  1001 => (x"33",x"54",x"41",x"46"),
  1002 => (x"20",x"20",x"20",x"32"),
  1003 => (x"00",x"00",x"00",x"00"),
  1004 => (x"31",x"54",x"41",x"46"),
  1005 => (x"20",x"20",x"20",x"36"),
  1006 => (x"d4",x"ff",x"1e",x"00"),
  1007 => (x"78",x"ff",x"c3",x"48"),
  1008 => (x"4f",x"26",x"48",x"68"),
  1009 => (x"48",x"d4",x"ff",x"1e"),
  1010 => (x"ff",x"78",x"ff",x"c3"),
  1011 => (x"e1",x"c0",x"48",x"d0"),
  1012 => (x"48",x"d4",x"ff",x"78"),
  1013 => (x"cb",x"c4",x"78",x"d4"),
  1014 => (x"d4",x"ff",x"48",x"e0"),
  1015 => (x"4f",x"26",x"50",x"bf"),
  1016 => (x"48",x"d0",x"ff",x"1e"),
  1017 => (x"26",x"78",x"e0",x"c0"),
  1018 => (x"cc",x"ff",x"1e",x"4f"),
  1019 => (x"99",x"49",x"70",x"87"),
  1020 => (x"c0",x"87",x"c6",x"02"),
  1021 => (x"f1",x"05",x"a9",x"fb"),
  1022 => (x"26",x"48",x"71",x"87"),
  1023 => (x"5b",x"5e",x"0e",x"4f"),
  1024 => (x"4b",x"71",x"0e",x"5c"),
  1025 => (x"f0",x"fe",x"4c",x"c0"),
  1026 => (x"99",x"49",x"70",x"87"),
  1027 => (x"87",x"f9",x"c0",x"02"),
  1028 => (x"02",x"a9",x"ec",x"c0"),
  1029 => (x"c0",x"87",x"f2",x"c0"),
  1030 => (x"c0",x"02",x"a9",x"fb"),
  1031 => (x"66",x"cc",x"87",x"eb"),
  1032 => (x"c7",x"03",x"ac",x"b7"),
  1033 => (x"02",x"66",x"d0",x"87"),
  1034 => (x"53",x"71",x"87",x"c2"),
  1035 => (x"c2",x"02",x"99",x"71"),
  1036 => (x"fe",x"84",x"c1",x"87"),
  1037 => (x"49",x"70",x"87",x"c3"),
  1038 => (x"87",x"cd",x"02",x"99"),
  1039 => (x"02",x"a9",x"ec",x"c0"),
  1040 => (x"fb",x"c0",x"87",x"c7"),
  1041 => (x"d5",x"ff",x"05",x"a9"),
  1042 => (x"02",x"66",x"d0",x"87"),
  1043 => (x"97",x"c0",x"87",x"c3"),
  1044 => (x"a9",x"ec",x"c0",x"7b"),
  1045 => (x"74",x"87",x"c4",x"05"),
  1046 => (x"74",x"87",x"c5",x"4a"),
  1047 => (x"8a",x"0a",x"c0",x"4a"),
  1048 => (x"4c",x"26",x"48",x"72"),
  1049 => (x"4f",x"26",x"4b",x"26"),
  1050 => (x"87",x"cd",x"fd",x"1e"),
  1051 => (x"c0",x"4a",x"49",x"70"),
  1052 => (x"c9",x"04",x"aa",x"f0"),
  1053 => (x"aa",x"f9",x"c0",x"87"),
  1054 => (x"c0",x"87",x"c3",x"01"),
  1055 => (x"c1",x"c1",x"8a",x"f0"),
  1056 => (x"87",x"c9",x"04",x"aa"),
  1057 => (x"01",x"aa",x"da",x"c1"),
  1058 => (x"f7",x"c0",x"87",x"c3"),
  1059 => (x"26",x"48",x"72",x"8a"),
  1060 => (x"5b",x"5e",x"0e",x"4f"),
  1061 => (x"4a",x"71",x"0e",x"5c"),
  1062 => (x"72",x"4c",x"d4",x"ff"),
  1063 => (x"87",x"ec",x"c0",x"49"),
  1064 => (x"02",x"9b",x"4b",x"70"),
  1065 => (x"8b",x"c1",x"87",x"c2"),
  1066 => (x"c5",x"48",x"d0",x"ff"),
  1067 => (x"7c",x"d5",x"c1",x"78"),
  1068 => (x"31",x"c6",x"49",x"73"),
  1069 => (x"97",x"dc",x"f2",x"c1"),
  1070 => (x"71",x"48",x"4a",x"bf"),
  1071 => (x"ff",x"7c",x"70",x"b0"),
  1072 => (x"78",x"c4",x"48",x"d0"),
  1073 => (x"4c",x"26",x"48",x"73"),
  1074 => (x"4f",x"26",x"4b",x"26"),
  1075 => (x"5c",x"5b",x"5e",x"0e"),
  1076 => (x"86",x"f8",x"0e",x"5d"),
  1077 => (x"a6",x"c4",x"4d",x"71"),
  1078 => (x"fb",x"78",x"c0",x"48"),
  1079 => (x"4b",x"c0",x"87",x"e6"),
  1080 => (x"97",x"cc",x"c6",x"c1"),
  1081 => (x"a9",x"c0",x"49",x"bf"),
  1082 => (x"fb",x"87",x"cf",x"04"),
  1083 => (x"83",x"c1",x"87",x"fb"),
  1084 => (x"97",x"cc",x"c6",x"c1"),
  1085 => (x"06",x"ab",x"49",x"bf"),
  1086 => (x"c6",x"c1",x"87",x"f1"),
  1087 => (x"02",x"bf",x"97",x"cc"),
  1088 => (x"f4",x"fa",x"87",x"cf"),
  1089 => (x"99",x"49",x"70",x"87"),
  1090 => (x"c0",x"87",x"c6",x"02"),
  1091 => (x"f1",x"05",x"a9",x"ec"),
  1092 => (x"75",x"4b",x"c0",x"87"),
  1093 => (x"87",x"e1",x"fa",x"7e"),
  1094 => (x"dc",x"fa",x"4c",x"70"),
  1095 => (x"fa",x"4d",x"70",x"87"),
  1096 => (x"4a",x"70",x"87",x"d7"),
  1097 => (x"49",x"6e",x"83",x"c1"),
  1098 => (x"69",x"97",x"81",x"c8"),
  1099 => (x"c7",x"02",x"ac",x"49"),
  1100 => (x"ac",x"ff",x"c0",x"87"),
  1101 => (x"87",x"e9",x"c0",x"05"),
  1102 => (x"81",x"c9",x"49",x"6e"),
  1103 => (x"ad",x"49",x"69",x"97"),
  1104 => (x"c0",x"87",x"c6",x"02"),
  1105 => (x"d8",x"05",x"ad",x"ff"),
  1106 => (x"ca",x"49",x"6e",x"87"),
  1107 => (x"49",x"69",x"97",x"81"),
  1108 => (x"87",x"c6",x"02",x"aa"),
  1109 => (x"05",x"aa",x"ff",x"c0"),
  1110 => (x"a6",x"c4",x"87",x"c7"),
  1111 => (x"d3",x"78",x"c1",x"48"),
  1112 => (x"ac",x"ec",x"c0",x"87"),
  1113 => (x"c0",x"87",x"c6",x"02"),
  1114 => (x"c7",x"05",x"ac",x"fb"),
  1115 => (x"c4",x"4b",x"c0",x"87"),
  1116 => (x"78",x"c1",x"48",x"a6"),
  1117 => (x"fe",x"02",x"66",x"c4"),
  1118 => (x"e3",x"f9",x"87",x"db"),
  1119 => (x"f8",x"48",x"73",x"87"),
  1120 => (x"26",x"4d",x"26",x"8e"),
  1121 => (x"26",x"4b",x"26",x"4c"),
  1122 => (x"00",x"00",x"00",x"4f"),
  1123 => (x"5b",x"5e",x"0e",x"00"),
  1124 => (x"f8",x"0e",x"5d",x"5c"),
  1125 => (x"ff",x"7e",x"71",x"86"),
  1126 => (x"1e",x"6e",x"4b",x"d4"),
  1127 => (x"49",x"e8",x"cb",x"c4"),
  1128 => (x"87",x"e3",x"df",x"ff"),
  1129 => (x"98",x"70",x"86",x"c4"),
  1130 => (x"87",x"d0",x"c4",x"02"),
  1131 => (x"c1",x"48",x"a6",x"c4"),
  1132 => (x"78",x"bf",x"e4",x"f2"),
  1133 => (x"d8",x"fb",x"49",x"6e"),
  1134 => (x"48",x"d0",x"ff",x"87"),
  1135 => (x"d6",x"c1",x"78",x"c5"),
  1136 => (x"6e",x"4a",x"c0",x"7b"),
  1137 => (x"11",x"81",x"72",x"49"),
  1138 => (x"cb",x"82",x"c1",x"7b"),
  1139 => (x"f2",x"04",x"aa",x"b7"),
  1140 => (x"c3",x"4a",x"cc",x"87"),
  1141 => (x"82",x"c1",x"7b",x"ff"),
  1142 => (x"aa",x"b7",x"e0",x"c0"),
  1143 => (x"ff",x"87",x"f4",x"04"),
  1144 => (x"78",x"c4",x"48",x"d0"),
  1145 => (x"c5",x"7b",x"ff",x"c3"),
  1146 => (x"7b",x"d3",x"c1",x"78"),
  1147 => (x"78",x"c4",x"7b",x"c1"),
  1148 => (x"66",x"c4",x"7e",x"73"),
  1149 => (x"a8",x"b7",x"c0",x"48"),
  1150 => (x"87",x"ee",x"c2",x"06"),
  1151 => (x"bf",x"f0",x"cb",x"c4"),
  1152 => (x"48",x"66",x"c4",x"4c"),
  1153 => (x"a6",x"c8",x"88",x"74"),
  1154 => (x"02",x"9c",x"74",x"58"),
  1155 => (x"c3",x"87",x"f7",x"c1"),
  1156 => (x"c8",x"4d",x"ec",x"fe"),
  1157 => (x"c0",x"8c",x"4b",x"c0"),
  1158 => (x"c6",x"03",x"ac",x"b7"),
  1159 => (x"a4",x"c0",x"c8",x"87"),
  1160 => (x"c4",x"4c",x"c0",x"4b"),
  1161 => (x"bf",x"97",x"e0",x"cb"),
  1162 => (x"02",x"99",x"d0",x"49"),
  1163 => (x"1e",x"c0",x"87",x"d1"),
  1164 => (x"49",x"e8",x"cb",x"c4"),
  1165 => (x"c4",x"87",x"d6",x"e2"),
  1166 => (x"4a",x"49",x"70",x"86"),
  1167 => (x"c3",x"87",x"eb",x"c0"),
  1168 => (x"c4",x"1e",x"ec",x"fe"),
  1169 => (x"e2",x"49",x"e8",x"cb"),
  1170 => (x"86",x"c4",x"87",x"c3"),
  1171 => (x"ff",x"4a",x"49",x"70"),
  1172 => (x"c5",x"c8",x"48",x"d0"),
  1173 => (x"c1",x"48",x"6e",x"78"),
  1174 => (x"48",x"15",x"78",x"d4"),
  1175 => (x"c1",x"78",x"08",x"6e"),
  1176 => (x"f5",x"ff",x"05",x"8b"),
  1177 => (x"48",x"d0",x"ff",x"87"),
  1178 => (x"9a",x"72",x"78",x"c4"),
  1179 => (x"c0",x"87",x"c5",x"05"),
  1180 => (x"87",x"ca",x"c1",x"48"),
  1181 => (x"cb",x"c4",x"1e",x"c1"),
  1182 => (x"df",x"ff",x"49",x"e8"),
  1183 => (x"86",x"c4",x"87",x"f0"),
  1184 => (x"fe",x"05",x"9c",x"74"),
  1185 => (x"66",x"c4",x"87",x"c9"),
  1186 => (x"a8",x"b7",x"c0",x"48"),
  1187 => (x"c4",x"87",x"d1",x"06"),
  1188 => (x"c0",x"48",x"e8",x"cb"),
  1189 => (x"c0",x"80",x"d0",x"78"),
  1190 => (x"c4",x"80",x"f4",x"78"),
  1191 => (x"78",x"bf",x"f4",x"cb"),
  1192 => (x"c0",x"48",x"66",x"c4"),
  1193 => (x"fd",x"01",x"a8",x"b7"),
  1194 => (x"4b",x"6e",x"87",x"d2"),
  1195 => (x"c5",x"48",x"d0",x"ff"),
  1196 => (x"7b",x"d3",x"c1",x"78"),
  1197 => (x"78",x"c4",x"7b",x"c0"),
  1198 => (x"87",x"c2",x"48",x"c1"),
  1199 => (x"8e",x"f8",x"48",x"c0"),
  1200 => (x"4c",x"26",x"4d",x"26"),
  1201 => (x"4f",x"26",x"4b",x"26"),
  1202 => (x"5c",x"5b",x"5e",x"0e"),
  1203 => (x"86",x"fc",x"0e",x"5d"),
  1204 => (x"4b",x"c0",x"4d",x"71"),
  1205 => (x"c0",x"04",x"ad",x"4c"),
  1206 => (x"c3",x"c1",x"87",x"e8"),
  1207 => (x"9c",x"74",x"1e",x"cc"),
  1208 => (x"c0",x"87",x"c4",x"02"),
  1209 => (x"c1",x"87",x"c2",x"4a"),
  1210 => (x"ea",x"49",x"72",x"4a"),
  1211 => (x"86",x"c4",x"87",x"ec"),
  1212 => (x"83",x"c1",x"7e",x"70"),
  1213 => (x"87",x"c2",x"05",x"6e"),
  1214 => (x"84",x"c1",x"4b",x"75"),
  1215 => (x"ff",x"06",x"ab",x"75"),
  1216 => (x"48",x"6e",x"87",x"d8"),
  1217 => (x"4d",x"26",x"8e",x"fc"),
  1218 => (x"4b",x"26",x"4c",x"26"),
  1219 => (x"71",x"1e",x"4f",x"26"),
  1220 => (x"ff",x"c3",x"49",x"4a"),
  1221 => (x"48",x"d4",x"ff",x"99"),
  1222 => (x"49",x"72",x"78",x"71"),
  1223 => (x"c3",x"29",x"b7",x"c8"),
  1224 => (x"78",x"71",x"99",x"ff"),
  1225 => (x"b7",x"d0",x"49",x"72"),
  1226 => (x"99",x"ff",x"c3",x"29"),
  1227 => (x"49",x"72",x"78",x"71"),
  1228 => (x"c3",x"29",x"b7",x"d8"),
  1229 => (x"78",x"71",x"99",x"ff"),
  1230 => (x"5e",x"0e",x"4f",x"26"),
  1231 => (x"0e",x"5d",x"5c",x"5b"),
  1232 => (x"4a",x"71",x"86",x"fc"),
  1233 => (x"49",x"72",x"4c",x"c0"),
  1234 => (x"87",x"ff",x"ec",x"c1"),
  1235 => (x"da",x"05",x"98",x"70"),
  1236 => (x"73",x"4b",x"c1",x"87"),
  1237 => (x"d2",x"ee",x"c1",x"49"),
  1238 => (x"05",x"98",x"70",x"87"),
  1239 => (x"4c",x"c1",x"87",x"c2"),
  1240 => (x"d1",x"c4",x"83",x"c1"),
  1241 => (x"ab",x"b7",x"bf",x"c4"),
  1242 => (x"ff",x"87",x"e8",x"06"),
  1243 => (x"e1",x"c8",x"48",x"d0"),
  1244 => (x"48",x"d4",x"ff",x"78"),
  1245 => (x"9c",x"74",x"78",x"dd"),
  1246 => (x"c4",x"87",x"c7",x"02"),
  1247 => (x"4d",x"bf",x"ec",x"d1"),
  1248 => (x"4d",x"c0",x"87",x"c2"),
  1249 => (x"c5",x"fe",x"49",x"75"),
  1250 => (x"02",x"9c",x"74",x"87"),
  1251 => (x"d1",x"c4",x"87",x"c7"),
  1252 => (x"c2",x"7e",x"bf",x"ec"),
  1253 => (x"6e",x"7e",x"c0",x"87"),
  1254 => (x"87",x"f2",x"fd",x"49"),
  1255 => (x"ed",x"fd",x"49",x"c0"),
  1256 => (x"fd",x"49",x"c0",x"87"),
  1257 => (x"d0",x"ff",x"87",x"e8"),
  1258 => (x"78",x"e0",x"c0",x"48"),
  1259 => (x"49",x"dc",x"1e",x"c1"),
  1260 => (x"87",x"da",x"fb",x"c0"),
  1261 => (x"8e",x"f8",x"48",x"74"),
  1262 => (x"4c",x"26",x"4d",x"26"),
  1263 => (x"4f",x"26",x"4b",x"26"),
  1264 => (x"c4",x"4a",x"71",x"1e"),
  1265 => (x"87",x"c9",x"02",x"66"),
  1266 => (x"89",x"c3",x"c1",x"49"),
  1267 => (x"cc",x"87",x"c9",x"02"),
  1268 => (x"f6",x"49",x"72",x"87"),
  1269 => (x"87",x"c5",x"87",x"f7"),
  1270 => (x"dd",x"fd",x"49",x"72"),
  1271 => (x"0e",x"4f",x"26",x"87"),
  1272 => (x"5d",x"5c",x"5b",x"5e"),
  1273 => (x"71",x"86",x"fc",x"0e"),
  1274 => (x"91",x"de",x"49",x"4c"),
  1275 => (x"4d",x"d0",x"cc",x"c4"),
  1276 => (x"6d",x"97",x"85",x"71"),
  1277 => (x"87",x"dc",x"c1",x"02"),
  1278 => (x"bf",x"fc",x"cb",x"c4"),
  1279 => (x"72",x"82",x"74",x"4a"),
  1280 => (x"87",x"c4",x"fb",x"49"),
  1281 => (x"02",x"6e",x"7e",x"70"),
  1282 => (x"c4",x"87",x"f2",x"c0"),
  1283 => (x"6e",x"4b",x"c4",x"cc"),
  1284 => (x"fe",x"49",x"cb",x"4a"),
  1285 => (x"74",x"87",x"e2",x"f2"),
  1286 => (x"c1",x"93",x"cc",x"4b"),
  1287 => (x"c4",x"83",x"f8",x"f2"),
  1288 => (x"e0",x"d1",x"c1",x"83"),
  1289 => (x"c1",x"49",x"74",x"7b"),
  1290 => (x"75",x"87",x"d1",x"cd"),
  1291 => (x"e0",x"f2",x"c1",x"7b"),
  1292 => (x"1e",x"49",x"bf",x"97"),
  1293 => (x"49",x"c4",x"cc",x"c4"),
  1294 => (x"c4",x"87",x"c5",x"fe"),
  1295 => (x"c1",x"49",x"74",x"86"),
  1296 => (x"c0",x"87",x"f9",x"cc"),
  1297 => (x"d4",x"ce",x"c1",x"49"),
  1298 => (x"e4",x"cb",x"c4",x"87"),
  1299 => (x"c1",x"78",x"c0",x"48"),
  1300 => (x"87",x"ef",x"dd",x"49"),
  1301 => (x"4d",x"26",x"8e",x"fc"),
  1302 => (x"4b",x"26",x"4c",x"26"),
  1303 => (x"00",x"00",x"4f",x"26"),
  1304 => (x"64",x"61",x"6f",x"4c"),
  1305 => (x"2e",x"67",x"6e",x"69"),
  1306 => (x"0e",x"00",x"2e",x"2e"),
  1307 => (x"0e",x"5c",x"5b",x"5e"),
  1308 => (x"c4",x"4a",x"4b",x"71"),
  1309 => (x"82",x"bf",x"fc",x"cb"),
  1310 => (x"cb",x"f9",x"49",x"72"),
  1311 => (x"9c",x"4c",x"70",x"87"),
  1312 => (x"49",x"87",x"c4",x"02"),
  1313 => (x"c4",x"87",x"d8",x"e3"),
  1314 => (x"c0",x"48",x"fc",x"cb"),
  1315 => (x"dc",x"49",x"c1",x"78"),
  1316 => (x"4c",x"26",x"87",x"f1"),
  1317 => (x"4f",x"26",x"4b",x"26"),
  1318 => (x"5c",x"5b",x"5e",x"0e"),
  1319 => (x"86",x"f4",x"0e",x"5d"),
  1320 => (x"4d",x"ec",x"fe",x"c3"),
  1321 => (x"a6",x"c4",x"4c",x"c0"),
  1322 => (x"c4",x"78",x"c0",x"48"),
  1323 => (x"49",x"bf",x"fc",x"cb"),
  1324 => (x"a9",x"c0",x"7e",x"75"),
  1325 => (x"87",x"fb",x"c0",x"06"),
  1326 => (x"fe",x"c3",x"7e",x"75"),
  1327 => (x"02",x"98",x"48",x"ec"),
  1328 => (x"c1",x"87",x"f0",x"c0"),
  1329 => (x"c8",x"1e",x"cc",x"c3"),
  1330 => (x"87",x"c4",x"02",x"66"),
  1331 => (x"87",x"c2",x"4d",x"c0"),
  1332 => (x"49",x"75",x"4d",x"c1"),
  1333 => (x"c4",x"87",x"c3",x"e3"),
  1334 => (x"c1",x"7e",x"70",x"86"),
  1335 => (x"48",x"66",x"c4",x"84"),
  1336 => (x"a6",x"c8",x"80",x"c1"),
  1337 => (x"fc",x"cb",x"c4",x"58"),
  1338 => (x"03",x"ac",x"49",x"bf"),
  1339 => (x"05",x"6e",x"87",x"c5"),
  1340 => (x"6e",x"87",x"d0",x"ff"),
  1341 => (x"75",x"4c",x"c0",x"4d"),
  1342 => (x"e0",x"c3",x"02",x"9d"),
  1343 => (x"cc",x"c3",x"c1",x"87"),
  1344 => (x"02",x"66",x"c8",x"1e"),
  1345 => (x"a6",x"cc",x"87",x"c7"),
  1346 => (x"c5",x"78",x"c0",x"48"),
  1347 => (x"48",x"a6",x"cc",x"87"),
  1348 => (x"66",x"cc",x"78",x"c1"),
  1349 => (x"87",x"c2",x"e2",x"49"),
  1350 => (x"7e",x"70",x"86",x"c4"),
  1351 => (x"e9",x"c2",x"02",x"6e"),
  1352 => (x"cb",x"49",x"6e",x"87"),
  1353 => (x"49",x"69",x"97",x"81"),
  1354 => (x"c1",x"02",x"99",x"d0"),
  1355 => (x"d1",x"c1",x"87",x"d6"),
  1356 => (x"49",x"74",x"4a",x"eb"),
  1357 => (x"f2",x"c1",x"91",x"cc"),
  1358 => (x"79",x"72",x"81",x"f8"),
  1359 => (x"ff",x"c3",x"81",x"c8"),
  1360 => (x"de",x"49",x"74",x"51"),
  1361 => (x"d0",x"cc",x"c4",x"91"),
  1362 => (x"c2",x"85",x"71",x"4d"),
  1363 => (x"c1",x"7d",x"97",x"c1"),
  1364 => (x"e0",x"c0",x"49",x"a5"),
  1365 => (x"fc",x"c6",x"c4",x"51"),
  1366 => (x"d2",x"02",x"bf",x"97"),
  1367 => (x"c2",x"84",x"c1",x"87"),
  1368 => (x"c6",x"c4",x"4b",x"a5"),
  1369 => (x"49",x"db",x"4a",x"fc"),
  1370 => (x"87",x"cd",x"ed",x"fe"),
  1371 => (x"cd",x"87",x"db",x"c1"),
  1372 => (x"51",x"c0",x"49",x"a5"),
  1373 => (x"a5",x"c2",x"84",x"c1"),
  1374 => (x"cb",x"4a",x"6e",x"4b"),
  1375 => (x"f8",x"ec",x"fe",x"49"),
  1376 => (x"87",x"c6",x"c1",x"87"),
  1377 => (x"4a",x"df",x"cf",x"c1"),
  1378 => (x"91",x"cc",x"49",x"74"),
  1379 => (x"81",x"f8",x"f2",x"c1"),
  1380 => (x"c6",x"c4",x"79",x"72"),
  1381 => (x"02",x"bf",x"97",x"fc"),
  1382 => (x"49",x"74",x"87",x"d8"),
  1383 => (x"84",x"c1",x"91",x"de"),
  1384 => (x"4b",x"d0",x"cc",x"c4"),
  1385 => (x"c6",x"c4",x"83",x"71"),
  1386 => (x"49",x"dd",x"4a",x"fc"),
  1387 => (x"87",x"c9",x"ec",x"fe"),
  1388 => (x"4b",x"74",x"87",x"d8"),
  1389 => (x"cc",x"c4",x"93",x"de"),
  1390 => (x"a3",x"cb",x"83",x"d0"),
  1391 => (x"c1",x"51",x"c0",x"49"),
  1392 => (x"4a",x"6e",x"73",x"84"),
  1393 => (x"eb",x"fe",x"49",x"cb"),
  1394 => (x"66",x"c4",x"87",x"ef"),
  1395 => (x"c8",x"80",x"c1",x"48"),
  1396 => (x"ac",x"c7",x"58",x"a6"),
  1397 => (x"87",x"c5",x"c0",x"03"),
  1398 => (x"e0",x"fc",x"05",x"6e"),
  1399 => (x"f4",x"48",x"74",x"87"),
  1400 => (x"26",x"4d",x"26",x"8e"),
  1401 => (x"26",x"4b",x"26",x"4c"),
  1402 => (x"1e",x"73",x"1e",x"4f"),
  1403 => (x"cc",x"49",x"4b",x"71"),
  1404 => (x"f8",x"f2",x"c1",x"91"),
  1405 => (x"4a",x"a1",x"c8",x"81"),
  1406 => (x"48",x"dc",x"f2",x"c1"),
  1407 => (x"a1",x"c9",x"50",x"12"),
  1408 => (x"cc",x"c6",x"c1",x"4a"),
  1409 => (x"ca",x"50",x"12",x"48"),
  1410 => (x"e0",x"f2",x"c1",x"81"),
  1411 => (x"c1",x"50",x"11",x"48"),
  1412 => (x"bf",x"97",x"e0",x"f2"),
  1413 => (x"49",x"c0",x"1e",x"49"),
  1414 => (x"c4",x"87",x"e5",x"f6"),
  1415 => (x"de",x"48",x"e4",x"cb"),
  1416 => (x"d6",x"49",x"c1",x"78"),
  1417 => (x"8e",x"fc",x"87",x"dd"),
  1418 => (x"4f",x"26",x"4b",x"26"),
  1419 => (x"49",x"4a",x"71",x"1e"),
  1420 => (x"f2",x"c1",x"91",x"cc"),
  1421 => (x"81",x"c8",x"81",x"f8"),
  1422 => (x"cb",x"c4",x"48",x"11"),
  1423 => (x"cb",x"c4",x"58",x"e8"),
  1424 => (x"78",x"c0",x"48",x"fc"),
  1425 => (x"fa",x"d5",x"49",x"c1"),
  1426 => (x"1e",x"4f",x"26",x"87"),
  1427 => (x"c6",x"c1",x"49",x"c0"),
  1428 => (x"4f",x"26",x"87",x"cb"),
  1429 => (x"02",x"99",x"71",x"1e"),
  1430 => (x"f4",x"c1",x"87",x"d2"),
  1431 => (x"50",x"c0",x"48",x"d4"),
  1432 => (x"d8",x"c1",x"80",x"f7"),
  1433 => (x"f2",x"c1",x"40",x"ec"),
  1434 => (x"87",x"ce",x"78",x"f0"),
  1435 => (x"48",x"d0",x"f4",x"c1"),
  1436 => (x"78",x"e8",x"f2",x"c1"),
  1437 => (x"d9",x"c1",x"80",x"fc"),
  1438 => (x"4f",x"26",x"78",x"cb"),
  1439 => (x"5c",x"5b",x"5e",x"0e"),
  1440 => (x"4a",x"4c",x"71",x"0e"),
  1441 => (x"f2",x"c1",x"92",x"cc"),
  1442 => (x"a2",x"c8",x"82",x"f8"),
  1443 => (x"4b",x"a2",x"c9",x"49"),
  1444 => (x"1e",x"4b",x"6b",x"97"),
  1445 => (x"1e",x"49",x"69",x"97"),
  1446 => (x"49",x"12",x"82",x"ca"),
  1447 => (x"87",x"ca",x"f1",x"c0"),
  1448 => (x"de",x"d4",x"49",x"c0"),
  1449 => (x"c1",x"49",x"74",x"87"),
  1450 => (x"f8",x"87",x"d1",x"c3"),
  1451 => (x"26",x"4c",x"26",x"8e"),
  1452 => (x"1e",x"4f",x"26",x"4b"),
  1453 => (x"4b",x"71",x"1e",x"73"),
  1454 => (x"87",x"c0",x"ff",x"49"),
  1455 => (x"fb",x"fe",x"49",x"73"),
  1456 => (x"26",x"4b",x"26",x"87"),
  1457 => (x"1e",x"73",x"1e",x"4f"),
  1458 => (x"a3",x"c6",x"4b",x"71"),
  1459 => (x"87",x"db",x"02",x"4a"),
  1460 => (x"d6",x"02",x"8a",x"c1"),
  1461 => (x"c1",x"02",x"8a",x"87"),
  1462 => (x"02",x"8a",x"87",x"da"),
  1463 => (x"8a",x"87",x"fc",x"c0"),
  1464 => (x"87",x"e1",x"c0",x"02"),
  1465 => (x"87",x"cb",x"02",x"8a"),
  1466 => (x"c7",x"87",x"db",x"c1"),
  1467 => (x"87",x"fc",x"fc",x"49"),
  1468 => (x"c4",x"87",x"de",x"c1"),
  1469 => (x"02",x"bf",x"fc",x"cb"),
  1470 => (x"48",x"87",x"cb",x"c1"),
  1471 => (x"cc",x"c4",x"88",x"c1"),
  1472 => (x"c1",x"c1",x"58",x"c0"),
  1473 => (x"c0",x"cc",x"c4",x"87"),
  1474 => (x"f9",x"c0",x"02",x"bf"),
  1475 => (x"fc",x"cb",x"c4",x"87"),
  1476 => (x"80",x"c1",x"48",x"bf"),
  1477 => (x"58",x"c0",x"cc",x"c4"),
  1478 => (x"c4",x"87",x"eb",x"c0"),
  1479 => (x"49",x"bf",x"fc",x"cb"),
  1480 => (x"cc",x"c4",x"89",x"c6"),
  1481 => (x"b7",x"c0",x"59",x"c0"),
  1482 => (x"87",x"da",x"03",x"a9"),
  1483 => (x"48",x"fc",x"cb",x"c4"),
  1484 => (x"87",x"d2",x"78",x"c0"),
  1485 => (x"bf",x"c0",x"cc",x"c4"),
  1486 => (x"c4",x"87",x"cb",x"02"),
  1487 => (x"48",x"bf",x"fc",x"cb"),
  1488 => (x"cc",x"c4",x"80",x"c6"),
  1489 => (x"49",x"c0",x"58",x"c0"),
  1490 => (x"73",x"87",x"f8",x"d1"),
  1491 => (x"eb",x"c0",x"c1",x"49"),
  1492 => (x"26",x"4b",x"26",x"87"),
  1493 => (x"5b",x"5e",x"0e",x"4f"),
  1494 => (x"ff",x"0e",x"5d",x"5c"),
  1495 => (x"a6",x"dc",x"86",x"d0"),
  1496 => (x"48",x"a6",x"c8",x"59"),
  1497 => (x"80",x"c4",x"78",x"c0"),
  1498 => (x"78",x"66",x"c4",x"c1"),
  1499 => (x"78",x"c1",x"80",x"c4"),
  1500 => (x"78",x"c1",x"80",x"c4"),
  1501 => (x"48",x"c0",x"cc",x"c4"),
  1502 => (x"cb",x"c4",x"78",x"c1"),
  1503 => (x"de",x"48",x"bf",x"e4"),
  1504 => (x"87",x"cb",x"05",x"a8"),
  1505 => (x"70",x"87",x"d1",x"f4"),
  1506 => (x"59",x"a6",x"cc",x"49"),
  1507 => (x"e0",x"87",x"ed",x"cf"),
  1508 => (x"d4",x"e1",x"87",x"f2"),
  1509 => (x"87",x"e1",x"e0",x"87"),
  1510 => (x"fb",x"c0",x"4c",x"70"),
  1511 => (x"f1",x"c1",x"02",x"ac"),
  1512 => (x"05",x"66",x"d8",x"87"),
  1513 => (x"c1",x"87",x"e2",x"c1"),
  1514 => (x"c4",x"4a",x"66",x"c0"),
  1515 => (x"c1",x"7e",x"6a",x"82"),
  1516 => (x"6e",x"48",x"f4",x"ee"),
  1517 => (x"20",x"41",x"20",x"49"),
  1518 => (x"c1",x"51",x"10",x"41"),
  1519 => (x"c1",x"48",x"66",x"c0"),
  1520 => (x"6a",x"78",x"e9",x"d7"),
  1521 => (x"74",x"81",x"c7",x"49"),
  1522 => (x"66",x"c0",x"c1",x"51"),
  1523 => (x"c1",x"81",x"c8",x"49"),
  1524 => (x"66",x"c0",x"c1",x"51"),
  1525 => (x"c0",x"81",x"c9",x"49"),
  1526 => (x"66",x"c0",x"c1",x"51"),
  1527 => (x"c0",x"81",x"ca",x"49"),
  1528 => (x"d8",x"1e",x"c1",x"51"),
  1529 => (x"c8",x"49",x"6a",x"1e"),
  1530 => (x"87",x"d1",x"e0",x"81"),
  1531 => (x"c4",x"c1",x"86",x"c8"),
  1532 => (x"a8",x"c0",x"48",x"66"),
  1533 => (x"c8",x"87",x"c7",x"01"),
  1534 => (x"78",x"c1",x"48",x"a6"),
  1535 => (x"c4",x"c1",x"87",x"cf"),
  1536 => (x"88",x"c1",x"48",x"66"),
  1537 => (x"c4",x"58",x"a6",x"d0"),
  1538 => (x"dc",x"df",x"ff",x"87"),
  1539 => (x"48",x"a6",x"d0",x"87"),
  1540 => (x"9c",x"74",x"78",x"c2"),
  1541 => (x"87",x"e0",x"cd",x"02"),
  1542 => (x"c1",x"48",x"66",x"c8"),
  1543 => (x"03",x"a8",x"66",x"c8"),
  1544 => (x"dc",x"87",x"d5",x"cd"),
  1545 => (x"78",x"c0",x"48",x"a6"),
  1546 => (x"cc",x"de",x"ff",x"7e"),
  1547 => (x"c1",x"4c",x"70",x"87"),
  1548 => (x"c2",x"05",x"ac",x"d0"),
  1549 => (x"a6",x"c4",x"87",x"da"),
  1550 => (x"e0",x"78",x"6e",x"48"),
  1551 => (x"49",x"70",x"87",x"ea"),
  1552 => (x"f4",x"dd",x"ff",x"7e"),
  1553 => (x"c0",x"4c",x"70",x"87"),
  1554 => (x"c1",x"05",x"ac",x"ec"),
  1555 => (x"66",x"c8",x"87",x"ed"),
  1556 => (x"c1",x"91",x"cc",x"49"),
  1557 => (x"c4",x"81",x"66",x"c0"),
  1558 => (x"4d",x"6a",x"4a",x"a1"),
  1559 => (x"6e",x"4a",x"a1",x"c8"),
  1560 => (x"ec",x"d8",x"c1",x"52"),
  1561 => (x"d0",x"dd",x"ff",x"79"),
  1562 => (x"9c",x"4c",x"70",x"87"),
  1563 => (x"c0",x"87",x"d9",x"02"),
  1564 => (x"d3",x"02",x"ac",x"fb"),
  1565 => (x"ff",x"55",x"74",x"87"),
  1566 => (x"70",x"87",x"fe",x"dc"),
  1567 => (x"c7",x"02",x"9c",x"4c"),
  1568 => (x"ac",x"fb",x"c0",x"87"),
  1569 => (x"87",x"ed",x"ff",x"05"),
  1570 => (x"c2",x"55",x"e0",x"c0"),
  1571 => (x"97",x"c0",x"55",x"c1"),
  1572 => (x"49",x"66",x"d8",x"7d"),
  1573 => (x"05",x"a9",x"66",x"c4"),
  1574 => (x"66",x"c8",x"87",x"db"),
  1575 => (x"a8",x"66",x"cc",x"48"),
  1576 => (x"c8",x"87",x"ca",x"04"),
  1577 => (x"80",x"c1",x"48",x"66"),
  1578 => (x"c8",x"58",x"a6",x"cc"),
  1579 => (x"48",x"66",x"cc",x"87"),
  1580 => (x"a6",x"d0",x"88",x"c1"),
  1581 => (x"c0",x"dc",x"ff",x"58"),
  1582 => (x"c1",x"4c",x"70",x"87"),
  1583 => (x"c8",x"05",x"ac",x"d0"),
  1584 => (x"48",x"66",x"d4",x"87"),
  1585 => (x"a6",x"d8",x"80",x"c1"),
  1586 => (x"ac",x"d0",x"c1",x"58"),
  1587 => (x"87",x"e6",x"fd",x"02"),
  1588 => (x"48",x"a6",x"e0",x"c0"),
  1589 => (x"6e",x"78",x"66",x"d8"),
  1590 => (x"66",x"e0",x"c0",x"48"),
  1591 => (x"e9",x"c9",x"05",x"a8"),
  1592 => (x"a6",x"e4",x"c0",x"87"),
  1593 => (x"e0",x"78",x"c0",x"48"),
  1594 => (x"74",x"78",x"c0",x"80"),
  1595 => (x"88",x"fb",x"c0",x"48"),
  1596 => (x"58",x"a6",x"ec",x"c0"),
  1597 => (x"c8",x"02",x"98",x"70"),
  1598 => (x"cb",x"48",x"87",x"ea"),
  1599 => (x"a6",x"ec",x"c0",x"88"),
  1600 => (x"02",x"98",x"70",x"58"),
  1601 => (x"48",x"87",x"d3",x"c1"),
  1602 => (x"ec",x"c0",x"88",x"c9"),
  1603 => (x"98",x"70",x"58",x"a6"),
  1604 => (x"87",x"ed",x"c3",x"02"),
  1605 => (x"c0",x"88",x"c4",x"48"),
  1606 => (x"70",x"58",x"a6",x"ec"),
  1607 => (x"87",x"d0",x"02",x"98"),
  1608 => (x"c0",x"88",x"c1",x"48"),
  1609 => (x"70",x"58",x"a6",x"ec"),
  1610 => (x"d4",x"c3",x"02",x"98"),
  1611 => (x"87",x"ee",x"c7",x"87"),
  1612 => (x"c0",x"48",x"a6",x"dc"),
  1613 => (x"d9",x"ff",x"78",x"f0"),
  1614 => (x"4c",x"70",x"87",x"ff"),
  1615 => (x"02",x"ac",x"ec",x"c0"),
  1616 => (x"c0",x"87",x"c4",x"c0"),
  1617 => (x"c0",x"5c",x"a6",x"e0"),
  1618 => (x"cd",x"02",x"ac",x"ec"),
  1619 => (x"e8",x"d9",x"ff",x"87"),
  1620 => (x"c0",x"4c",x"70",x"87"),
  1621 => (x"ff",x"05",x"ac",x"ec"),
  1622 => (x"ec",x"c0",x"87",x"f3"),
  1623 => (x"c4",x"c0",x"02",x"ac"),
  1624 => (x"d4",x"d9",x"ff",x"87"),
  1625 => (x"ca",x"1e",x"c0",x"87"),
  1626 => (x"49",x"66",x"d0",x"1e"),
  1627 => (x"c8",x"c1",x"91",x"cc"),
  1628 => (x"80",x"71",x"48",x"66"),
  1629 => (x"c8",x"58",x"a6",x"cc"),
  1630 => (x"80",x"c4",x"48",x"66"),
  1631 => (x"cc",x"58",x"a6",x"d0"),
  1632 => (x"ff",x"49",x"bf",x"66"),
  1633 => (x"c1",x"87",x"f6",x"d9"),
  1634 => (x"d4",x"1e",x"de",x"1e"),
  1635 => (x"ff",x"49",x"bf",x"66"),
  1636 => (x"d0",x"87",x"ea",x"d9"),
  1637 => (x"c0",x"49",x"70",x"86"),
  1638 => (x"ec",x"c0",x"89",x"09"),
  1639 => (x"e8",x"c0",x"59",x"a6"),
  1640 => (x"a8",x"c0",x"48",x"66"),
  1641 => (x"87",x"ee",x"c0",x"06"),
  1642 => (x"48",x"66",x"e8",x"c0"),
  1643 => (x"c0",x"03",x"a8",x"dd"),
  1644 => (x"66",x"c4",x"87",x"e4"),
  1645 => (x"e8",x"c0",x"49",x"bf"),
  1646 => (x"e0",x"c0",x"81",x"66"),
  1647 => (x"66",x"e8",x"c0",x"51"),
  1648 => (x"c4",x"81",x"c1",x"49"),
  1649 => (x"c2",x"81",x"bf",x"66"),
  1650 => (x"e8",x"c0",x"51",x"c1"),
  1651 => (x"81",x"c2",x"49",x"66"),
  1652 => (x"81",x"bf",x"66",x"c4"),
  1653 => (x"48",x"6e",x"51",x"c0"),
  1654 => (x"78",x"e9",x"d7",x"c1"),
  1655 => (x"81",x"c8",x"49",x"6e"),
  1656 => (x"6e",x"51",x"66",x"d0"),
  1657 => (x"d4",x"81",x"c9",x"49"),
  1658 => (x"49",x"6e",x"51",x"66"),
  1659 => (x"66",x"dc",x"81",x"ca"),
  1660 => (x"48",x"66",x"d0",x"51"),
  1661 => (x"a6",x"d4",x"80",x"c1"),
  1662 => (x"80",x"f4",x"48",x"58"),
  1663 => (x"e3",x"c4",x"78",x"c1"),
  1664 => (x"e3",x"d9",x"ff",x"87"),
  1665 => (x"c0",x"49",x"70",x"87"),
  1666 => (x"ff",x"59",x"a6",x"ec"),
  1667 => (x"70",x"87",x"d9",x"d9"),
  1668 => (x"a6",x"e0",x"c0",x"49"),
  1669 => (x"48",x"66",x"dc",x"59"),
  1670 => (x"05",x"a8",x"ec",x"c0"),
  1671 => (x"dc",x"87",x"ca",x"c0"),
  1672 => (x"e8",x"c0",x"48",x"a6"),
  1673 => (x"c4",x"c0",x"78",x"66"),
  1674 => (x"cc",x"d6",x"ff",x"87"),
  1675 => (x"49",x"66",x"c8",x"87"),
  1676 => (x"c0",x"c1",x"91",x"cc"),
  1677 => (x"80",x"71",x"48",x"66"),
  1678 => (x"c4",x"58",x"a6",x"c8"),
  1679 => (x"82",x"c8",x"4a",x"66"),
  1680 => (x"ca",x"49",x"66",x"c4"),
  1681 => (x"66",x"e8",x"c0",x"81"),
  1682 => (x"49",x"66",x"dc",x"51"),
  1683 => (x"e8",x"c0",x"81",x"c1"),
  1684 => (x"48",x"c1",x"89",x"66"),
  1685 => (x"49",x"70",x"30",x"71"),
  1686 => (x"97",x"71",x"89",x"c1"),
  1687 => (x"d4",x"d0",x"c4",x"7a"),
  1688 => (x"e8",x"c0",x"49",x"bf"),
  1689 => (x"6a",x"97",x"29",x"66"),
  1690 => (x"98",x"71",x"48",x"4a"),
  1691 => (x"58",x"a6",x"f0",x"c0"),
  1692 => (x"c4",x"49",x"66",x"c4"),
  1693 => (x"c0",x"4d",x"69",x"81"),
  1694 => (x"6e",x"48",x"66",x"e0"),
  1695 => (x"c5",x"c0",x"02",x"a8"),
  1696 => (x"c0",x"7e",x"c0",x"87"),
  1697 => (x"7e",x"c1",x"87",x"c2"),
  1698 => (x"e0",x"c0",x"1e",x"6e"),
  1699 => (x"ff",x"49",x"75",x"1e"),
  1700 => (x"c8",x"87",x"ea",x"d5"),
  1701 => (x"c0",x"4c",x"70",x"86"),
  1702 => (x"c1",x"06",x"ac",x"b7"),
  1703 => (x"85",x"74",x"87",x"d0"),
  1704 => (x"74",x"49",x"e0",x"c0"),
  1705 => (x"c1",x"4b",x"75",x"89"),
  1706 => (x"71",x"4a",x"c0",x"ef"),
  1707 => (x"87",x"c9",x"d8",x"fe"),
  1708 => (x"7e",x"75",x"85",x"c2"),
  1709 => (x"48",x"66",x"e4",x"c0"),
  1710 => (x"e8",x"c0",x"80",x"c1"),
  1711 => (x"ec",x"c0",x"58",x"a6"),
  1712 => (x"81",x"c1",x"49",x"66"),
  1713 => (x"c0",x"02",x"a9",x"70"),
  1714 => (x"4d",x"c0",x"87",x"c5"),
  1715 => (x"c1",x"87",x"c2",x"c0"),
  1716 => (x"c2",x"1e",x"75",x"4d"),
  1717 => (x"e0",x"c0",x"49",x"a4"),
  1718 => (x"70",x"88",x"71",x"48"),
  1719 => (x"66",x"c8",x"1e",x"49"),
  1720 => (x"d8",x"d4",x"ff",x"49"),
  1721 => (x"c0",x"86",x"c8",x"87"),
  1722 => (x"ff",x"01",x"a8",x"b7"),
  1723 => (x"e4",x"c0",x"87",x"c6"),
  1724 => (x"d3",x"c0",x"02",x"66"),
  1725 => (x"49",x"66",x"c4",x"87"),
  1726 => (x"e4",x"c0",x"81",x"c9"),
  1727 => (x"66",x"c4",x"51",x"66"),
  1728 => (x"fc",x"d9",x"c1",x"48"),
  1729 => (x"87",x"ce",x"c0",x"78"),
  1730 => (x"c9",x"49",x"66",x"c4"),
  1731 => (x"c4",x"51",x"c2",x"81"),
  1732 => (x"da",x"c1",x"48",x"66"),
  1733 => (x"a6",x"c4",x"78",x"f3"),
  1734 => (x"c0",x"78",x"c1",x"48"),
  1735 => (x"d3",x"ff",x"87",x"c6"),
  1736 => (x"4c",x"70",x"87",x"c7"),
  1737 => (x"c0",x"02",x"66",x"c4"),
  1738 => (x"66",x"c8",x"87",x"f5"),
  1739 => (x"a8",x"66",x"cc",x"48"),
  1740 => (x"87",x"cb",x"c0",x"04"),
  1741 => (x"c1",x"48",x"66",x"c8"),
  1742 => (x"58",x"a6",x"cc",x"80"),
  1743 => (x"cc",x"87",x"e0",x"c0"),
  1744 => (x"88",x"c1",x"48",x"66"),
  1745 => (x"c0",x"58",x"a6",x"d0"),
  1746 => (x"c6",x"c1",x"87",x"d5"),
  1747 => (x"c8",x"c0",x"05",x"ac"),
  1748 => (x"48",x"66",x"d0",x"87"),
  1749 => (x"a6",x"d4",x"80",x"c1"),
  1750 => (x"cc",x"d2",x"ff",x"58"),
  1751 => (x"d4",x"4c",x"70",x"87"),
  1752 => (x"80",x"c1",x"48",x"66"),
  1753 => (x"74",x"58",x"a6",x"d8"),
  1754 => (x"cb",x"c0",x"02",x"9c"),
  1755 => (x"48",x"66",x"c8",x"87"),
  1756 => (x"a8",x"66",x"c8",x"c1"),
  1757 => (x"87",x"eb",x"f2",x"04"),
  1758 => (x"87",x"e4",x"d1",x"ff"),
  1759 => (x"c7",x"48",x"66",x"c8"),
  1760 => (x"e1",x"c0",x"03",x"a8"),
  1761 => (x"4c",x"66",x"c8",x"87"),
  1762 => (x"48",x"c0",x"cc",x"c4"),
  1763 => (x"49",x"74",x"78",x"c0"),
  1764 => (x"c0",x"c1",x"91",x"cc"),
  1765 => (x"a1",x"c4",x"81",x"66"),
  1766 => (x"c0",x"4a",x"6a",x"4a"),
  1767 => (x"84",x"c1",x"79",x"52"),
  1768 => (x"ff",x"04",x"ac",x"c7"),
  1769 => (x"d0",x"ff",x"87",x"e2"),
  1770 => (x"26",x"4d",x"26",x"8e"),
  1771 => (x"26",x"4b",x"26",x"4c"),
  1772 => (x"00",x"00",x"00",x"4f"),
  1773 => (x"64",x"61",x"6f",x"4c"),
  1774 => (x"20",x"2e",x"2a",x"20"),
  1775 => (x"00",x"00",x"00",x"00"),
  1776 => (x"1e",x"00",x"20",x"3a"),
  1777 => (x"4b",x"71",x"1e",x"73"),
  1778 => (x"87",x"c6",x"02",x"9b"),
  1779 => (x"48",x"fc",x"cb",x"c4"),
  1780 => (x"1e",x"c7",x"78",x"c0"),
  1781 => (x"bf",x"fc",x"cb",x"c4"),
  1782 => (x"f2",x"c1",x"1e",x"49"),
  1783 => (x"cb",x"c4",x"1e",x"f8"),
  1784 => (x"ed",x"49",x"bf",x"e4"),
  1785 => (x"86",x"cc",x"87",x"ef"),
  1786 => (x"bf",x"e4",x"cb",x"c4"),
  1787 => (x"87",x"e4",x"e9",x"49"),
  1788 => (x"c8",x"02",x"9b",x"73"),
  1789 => (x"f8",x"f2",x"c1",x"87"),
  1790 => (x"cd",x"ef",x"c0",x"49"),
  1791 => (x"26",x"4b",x"26",x"87"),
  1792 => (x"ec",x"cc",x"1e",x"4f"),
  1793 => (x"fe",x"49",x"c1",x"87"),
  1794 => (x"e2",x"fe",x"87",x"f9"),
  1795 => (x"98",x"70",x"87",x"d7"),
  1796 => (x"fe",x"87",x"cd",x"02"),
  1797 => (x"70",x"87",x"fe",x"e9"),
  1798 => (x"87",x"c4",x"02",x"98"),
  1799 => (x"87",x"c2",x"4a",x"c1"),
  1800 => (x"9a",x"72",x"4a",x"c0"),
  1801 => (x"c0",x"87",x"ce",x"05"),
  1802 => (x"d8",x"f1",x"c1",x"1e"),
  1803 => (x"d1",x"fc",x"c0",x"49"),
  1804 => (x"fe",x"86",x"c4",x"87"),
  1805 => (x"e5",x"cb",x"c2",x"87"),
  1806 => (x"c1",x"1e",x"c0",x"87"),
  1807 => (x"c0",x"49",x"e4",x"f1"),
  1808 => (x"c0",x"87",x"ff",x"fb"),
  1809 => (x"ff",x"cb",x"c2",x"1e"),
  1810 => (x"c0",x"49",x"70",x"87"),
  1811 => (x"c3",x"87",x"f3",x"fb"),
  1812 => (x"8e",x"f8",x"87",x"ea"),
  1813 => (x"00",x"00",x"4f",x"26"),
  1814 => (x"66",x"20",x"44",x"53"),
  1815 => (x"65",x"6c",x"69",x"61"),
  1816 => (x"00",x"00",x"2e",x"64"),
  1817 => (x"74",x"6f",x"6f",x"42"),
  1818 => (x"2e",x"67",x"6e",x"69"),
  1819 => (x"1e",x"00",x"2e",x"2e"),
  1820 => (x"e7",x"d0",x"49",x"c0"),
  1821 => (x"ed",x"c6",x"c2",x"87"),
  1822 => (x"f6",x"f1",x"c0",x"87"),
  1823 => (x"e5",x"c6",x"c2",x"87"),
  1824 => (x"26",x"87",x"ed",x"87"),
  1825 => (x"cb",x"c4",x"1e",x"4f"),
  1826 => (x"78",x"c0",x"48",x"fc"),
  1827 => (x"48",x"e4",x"cb",x"c4"),
  1828 => (x"ec",x"fd",x"78",x"c0"),
  1829 => (x"87",x"d7",x"ff",x"87"),
  1830 => (x"4f",x"26",x"48",x"c0"),
  1831 => (x"00",x"00",x"00",x"00"),
  1832 => (x"00",x"00",x"00",x"00"),
  1833 => (x"00",x"00",x"00",x"01"),
  1834 => (x"78",x"45",x"20",x"80"),
  1835 => (x"00",x"00",x"74",x"69"),
  1836 => (x"61",x"42",x"20",x"80"),
  1837 => (x"00",x"00",x"6b",x"63"),
  1838 => (x"00",x"00",x"16",x"2c"),
  1839 => (x"00",x"00",x"43",x"10"),
  1840 => (x"00",x"00",x"00",x"00"),
  1841 => (x"00",x"00",x"16",x"2c"),
  1842 => (x"00",x"00",x"43",x"2e"),
  1843 => (x"00",x"00",x"00",x"00"),
  1844 => (x"00",x"00",x"16",x"2c"),
  1845 => (x"00",x"00",x"43",x"4c"),
  1846 => (x"00",x"00",x"00",x"00"),
  1847 => (x"00",x"00",x"16",x"2c"),
  1848 => (x"00",x"00",x"43",x"6a"),
  1849 => (x"00",x"00",x"00",x"00"),
  1850 => (x"00",x"00",x"16",x"2c"),
  1851 => (x"00",x"00",x"43",x"88"),
  1852 => (x"00",x"00",x"00",x"00"),
  1853 => (x"00",x"00",x"16",x"2c"),
  1854 => (x"00",x"00",x"43",x"a6"),
  1855 => (x"00",x"00",x"00",x"00"),
  1856 => (x"00",x"00",x"16",x"2c"),
  1857 => (x"00",x"00",x"43",x"c4"),
  1858 => (x"00",x"00",x"00",x"00"),
  1859 => (x"00",x"00",x"16",x"2c"),
  1860 => (x"00",x"00",x"00",x"00"),
  1861 => (x"00",x"00",x"00",x"00"),
  1862 => (x"00",x"00",x"16",x"c5"),
  1863 => (x"00",x"00",x"00",x"00"),
  1864 => (x"00",x"00",x"00",x"00"),
  1865 => (x"48",x"f0",x"fe",x"1e"),
  1866 => (x"09",x"cd",x"78",x"c0"),
  1867 => (x"4f",x"26",x"09",x"79"),
  1868 => (x"fe",x"86",x"fc",x"1e"),
  1869 => (x"48",x"7e",x"bf",x"f0"),
  1870 => (x"4f",x"26",x"8e",x"fc"),
  1871 => (x"48",x"f0",x"fe",x"1e"),
  1872 => (x"4f",x"26",x"78",x"c1"),
  1873 => (x"48",x"f0",x"fe",x"1e"),
  1874 => (x"4f",x"26",x"78",x"c0"),
  1875 => (x"c0",x"4a",x"71",x"1e"),
  1876 => (x"a2",x"c1",x"7a",x"97"),
  1877 => (x"ca",x"51",x"c0",x"49"),
  1878 => (x"51",x"c0",x"49",x"a2"),
  1879 => (x"c0",x"49",x"a2",x"cb"),
  1880 => (x"0e",x"4f",x"26",x"51"),
  1881 => (x"0e",x"5c",x"5b",x"5e"),
  1882 => (x"4c",x"71",x"86",x"f0"),
  1883 => (x"97",x"49",x"a4",x"ca"),
  1884 => (x"a4",x"cb",x"7e",x"69"),
  1885 => (x"48",x"6b",x"97",x"4b"),
  1886 => (x"c1",x"58",x"a6",x"c8"),
  1887 => (x"58",x"a6",x"cc",x"80"),
  1888 => (x"a6",x"d0",x"98",x"c7"),
  1889 => (x"cc",x"48",x"6e",x"58"),
  1890 => (x"db",x"05",x"a8",x"66"),
  1891 => (x"7e",x"69",x"97",x"87"),
  1892 => (x"c8",x"48",x"6b",x"97"),
  1893 => (x"80",x"c1",x"58",x"a6"),
  1894 => (x"c7",x"58",x"a6",x"cc"),
  1895 => (x"58",x"a6",x"d0",x"98"),
  1896 => (x"66",x"cc",x"48",x"6e"),
  1897 => (x"87",x"e5",x"02",x"a8"),
  1898 => (x"cc",x"87",x"d9",x"fe"),
  1899 => (x"6b",x"97",x"4a",x"a4"),
  1900 => (x"49",x"a1",x"72",x"49"),
  1901 => (x"97",x"51",x"66",x"dc"),
  1902 => (x"48",x"6e",x"7e",x"6b"),
  1903 => (x"a6",x"c8",x"80",x"c1"),
  1904 => (x"cc",x"98",x"c7",x"58"),
  1905 => (x"97",x"70",x"58",x"a6"),
  1906 => (x"87",x"d1",x"c2",x"7b"),
  1907 => (x"f0",x"87",x"ed",x"fd"),
  1908 => (x"26",x"4c",x"26",x"8e"),
  1909 => (x"0e",x"4f",x"26",x"4b"),
  1910 => (x"5d",x"5c",x"5b",x"5e"),
  1911 => (x"71",x"86",x"f4",x"0e"),
  1912 => (x"7e",x"6d",x"97",x"4d"),
  1913 => (x"97",x"4c",x"a5",x"c1"),
  1914 => (x"a6",x"c8",x"48",x"6c"),
  1915 => (x"c4",x"48",x"6e",x"58"),
  1916 => (x"c5",x"05",x"a8",x"66"),
  1917 => (x"c0",x"48",x"ff",x"87"),
  1918 => (x"c7",x"fd",x"87",x"e6"),
  1919 => (x"49",x"a5",x"c2",x"87"),
  1920 => (x"71",x"4b",x"6c",x"97"),
  1921 => (x"6b",x"97",x"4b",x"a3"),
  1922 => (x"7e",x"6c",x"97",x"4b"),
  1923 => (x"80",x"c1",x"48",x"6e"),
  1924 => (x"c7",x"58",x"a6",x"c8"),
  1925 => (x"58",x"a6",x"cc",x"98"),
  1926 => (x"fc",x"7c",x"97",x"70"),
  1927 => (x"48",x"73",x"87",x"de"),
  1928 => (x"4d",x"26",x"8e",x"f4"),
  1929 => (x"4b",x"26",x"4c",x"26"),
  1930 => (x"5e",x"0e",x"4f",x"26"),
  1931 => (x"f4",x"0e",x"5c",x"5b"),
  1932 => (x"d8",x"4c",x"71",x"86"),
  1933 => (x"ff",x"c3",x"4a",x"66"),
  1934 => (x"4b",x"a4",x"c2",x"9a"),
  1935 => (x"73",x"49",x"6c",x"97"),
  1936 => (x"51",x"72",x"49",x"a1"),
  1937 => (x"6e",x"7e",x"6c",x"97"),
  1938 => (x"c8",x"80",x"c1",x"48"),
  1939 => (x"98",x"c7",x"58",x"a6"),
  1940 => (x"70",x"58",x"a6",x"cc"),
  1941 => (x"26",x"8e",x"f4",x"54"),
  1942 => (x"26",x"4b",x"26",x"4c"),
  1943 => (x"1e",x"73",x"1e",x"4f"),
  1944 => (x"df",x"fb",x"86",x"f4"),
  1945 => (x"4b",x"bf",x"e0",x"87"),
  1946 => (x"c0",x"e0",x"c0",x"49"),
  1947 => (x"87",x"cb",x"02",x"99"),
  1948 => (x"cf",x"c4",x"1e",x"73"),
  1949 => (x"f1",x"fe",x"49",x"e4"),
  1950 => (x"73",x"86",x"c4",x"87"),
  1951 => (x"99",x"c0",x"d0",x"49"),
  1952 => (x"87",x"c0",x"c1",x"02"),
  1953 => (x"97",x"ee",x"cf",x"c4"),
  1954 => (x"cf",x"c4",x"7e",x"bf"),
  1955 => (x"48",x"bf",x"97",x"ef"),
  1956 => (x"6e",x"58",x"a6",x"c8"),
  1957 => (x"a8",x"66",x"c4",x"48"),
  1958 => (x"87",x"e8",x"c0",x"02"),
  1959 => (x"97",x"ee",x"cf",x"c4"),
  1960 => (x"cf",x"c4",x"49",x"bf"),
  1961 => (x"48",x"11",x"81",x"f0"),
  1962 => (x"c4",x"78",x"08",x"e0"),
  1963 => (x"bf",x"97",x"ee",x"cf"),
  1964 => (x"c1",x"48",x"6e",x"7e"),
  1965 => (x"58",x"a6",x"c8",x"80"),
  1966 => (x"a6",x"cc",x"98",x"c7"),
  1967 => (x"ee",x"cf",x"c4",x"58"),
  1968 => (x"50",x"66",x"c8",x"48"),
  1969 => (x"49",x"4b",x"bf",x"e4"),
  1970 => (x"99",x"c0",x"e0",x"c0"),
  1971 => (x"73",x"87",x"cb",x"02"),
  1972 => (x"f8",x"cf",x"c4",x"1e"),
  1973 => (x"87",x"d2",x"fd",x"49"),
  1974 => (x"49",x"73",x"86",x"c4"),
  1975 => (x"02",x"99",x"c0",x"d0"),
  1976 => (x"c4",x"87",x"c0",x"c1"),
  1977 => (x"bf",x"97",x"c2",x"d0"),
  1978 => (x"c3",x"d0",x"c4",x"7e"),
  1979 => (x"c8",x"48",x"bf",x"97"),
  1980 => (x"48",x"6e",x"58",x"a6"),
  1981 => (x"02",x"a8",x"66",x"c4"),
  1982 => (x"c4",x"87",x"e8",x"c0"),
  1983 => (x"bf",x"97",x"c2",x"d0"),
  1984 => (x"c4",x"d0",x"c4",x"49"),
  1985 => (x"e4",x"48",x"11",x"81"),
  1986 => (x"d0",x"c4",x"78",x"08"),
  1987 => (x"7e",x"bf",x"97",x"c2"),
  1988 => (x"80",x"c1",x"48",x"6e"),
  1989 => (x"c7",x"58",x"a6",x"c8"),
  1990 => (x"58",x"a6",x"cc",x"98"),
  1991 => (x"48",x"c2",x"d0",x"c4"),
  1992 => (x"f8",x"50",x"66",x"c8"),
  1993 => (x"7e",x"70",x"87",x"ca"),
  1994 => (x"f4",x"87",x"d1",x"f8"),
  1995 => (x"26",x"4b",x"26",x"8e"),
  1996 => (x"cf",x"c4",x"1e",x"4f"),
  1997 => (x"d3",x"f8",x"49",x"e4"),
  1998 => (x"f8",x"cf",x"c4",x"87"),
  1999 => (x"87",x"cc",x"f8",x"49"),
  2000 => (x"49",x"dd",x"f9",x"c1"),
  2001 => (x"c2",x"87",x"dd",x"f7"),
  2002 => (x"4f",x"26",x"87",x"fb"),
  2003 => (x"c4",x"1e",x"73",x"1e"),
  2004 => (x"fa",x"49",x"e4",x"cf"),
  2005 => (x"4a",x"70",x"87",x"c1"),
  2006 => (x"04",x"aa",x"b7",x"c0"),
  2007 => (x"c3",x"87",x"cc",x"c2"),
  2008 => (x"c9",x"05",x"aa",x"f0"),
  2009 => (x"f4",x"ff",x"c1",x"87"),
  2010 => (x"c1",x"78",x"c1",x"48"),
  2011 => (x"e0",x"c3",x"87",x"ed"),
  2012 => (x"87",x"c9",x"05",x"aa"),
  2013 => (x"48",x"f8",x"ff",x"c1"),
  2014 => (x"de",x"c1",x"78",x"c1"),
  2015 => (x"f8",x"ff",x"c1",x"87"),
  2016 => (x"87",x"c6",x"02",x"bf"),
  2017 => (x"4b",x"a2",x"c0",x"c2"),
  2018 => (x"4b",x"72",x"87",x"c2"),
  2019 => (x"bf",x"f4",x"ff",x"c1"),
  2020 => (x"87",x"e0",x"c0",x"02"),
  2021 => (x"b7",x"c4",x"49",x"73"),
  2022 => (x"c1",x"c2",x"91",x"29"),
  2023 => (x"4a",x"73",x"81",x"dc"),
  2024 => (x"92",x"c2",x"9a",x"cf"),
  2025 => (x"30",x"72",x"48",x"c1"),
  2026 => (x"ba",x"ff",x"4a",x"70"),
  2027 => (x"98",x"69",x"48",x"72"),
  2028 => (x"87",x"db",x"79",x"70"),
  2029 => (x"b7",x"c4",x"49",x"73"),
  2030 => (x"c1",x"c2",x"91",x"29"),
  2031 => (x"4a",x"73",x"81",x"dc"),
  2032 => (x"92",x"c2",x"9a",x"cf"),
  2033 => (x"30",x"72",x"48",x"c3"),
  2034 => (x"69",x"48",x"4a",x"70"),
  2035 => (x"c1",x"79",x"70",x"b0"),
  2036 => (x"c0",x"48",x"f8",x"ff"),
  2037 => (x"f4",x"ff",x"c1",x"78"),
  2038 => (x"c4",x"78",x"c0",x"48"),
  2039 => (x"f7",x"49",x"e4",x"cf"),
  2040 => (x"4a",x"70",x"87",x"f5"),
  2041 => (x"03",x"aa",x"b7",x"c0"),
  2042 => (x"c0",x"87",x"f4",x"fd"),
  2043 => (x"26",x"4b",x"26",x"48"),
  2044 => (x"00",x"00",x"00",x"4f"),
  2045 => (x"00",x"00",x"00",x"00"),
  2046 => (x"00",x"00",x"00",x"00"),
  2047 => (x"49",x"4a",x"71",x"1e"),
  2048 => (x"26",x"87",x"c9",x"fd"),
  2049 => (x"4a",x"c0",x"1e",x"4f"),
  2050 => (x"91",x"c4",x"49",x"72"),
  2051 => (x"81",x"dc",x"c1",x"c2"),
  2052 => (x"82",x"c1",x"79",x"c0"),
  2053 => (x"04",x"aa",x"b7",x"d0"),
  2054 => (x"4f",x"26",x"87",x"ee"),
  2055 => (x"5c",x"5b",x"5e",x"0e"),
  2056 => (x"4d",x"71",x"0e",x"5d"),
  2057 => (x"75",x"87",x"dd",x"f4"),
  2058 => (x"2a",x"b7",x"c4",x"4a"),
  2059 => (x"dc",x"c1",x"c2",x"92"),
  2060 => (x"cf",x"4c",x"75",x"82"),
  2061 => (x"6a",x"94",x"c2",x"9c"),
  2062 => (x"2b",x"74",x"4b",x"49"),
  2063 => (x"48",x"c2",x"9b",x"c3"),
  2064 => (x"4c",x"70",x"30",x"74"),
  2065 => (x"48",x"74",x"bc",x"ff"),
  2066 => (x"7a",x"70",x"98",x"71"),
  2067 => (x"73",x"87",x"ed",x"f3"),
  2068 => (x"26",x"4d",x"26",x"48"),
  2069 => (x"26",x"4b",x"26",x"4c"),
  2070 => (x"00",x"00",x"00",x"4f"),
  2071 => (x"00",x"00",x"00",x"00"),
  2072 => (x"00",x"00",x"00",x"00"),
  2073 => (x"00",x"00",x"00",x"00"),
  2074 => (x"00",x"00",x"00",x"00"),
  2075 => (x"00",x"00",x"00",x"00"),
  2076 => (x"00",x"00",x"00",x"00"),
  2077 => (x"00",x"00",x"00",x"00"),
  2078 => (x"00",x"00",x"00",x"00"),
  2079 => (x"00",x"00",x"00",x"00"),
  2080 => (x"00",x"00",x"00",x"00"),
  2081 => (x"00",x"00",x"00",x"00"),
  2082 => (x"00",x"00",x"00",x"00"),
  2083 => (x"00",x"00",x"00",x"00"),
  2084 => (x"00",x"00",x"00",x"00"),
  2085 => (x"00",x"00",x"00",x"00"),
  2086 => (x"00",x"00",x"00",x"00"),
  2087 => (x"5c",x"5b",x"5e",x"0e"),
  2088 => (x"4a",x"71",x"0e",x"5d"),
  2089 => (x"72",x"4d",x"d4",x"ff"),
  2090 => (x"87",x"c6",x"02",x"9a"),
  2091 => (x"48",x"d8",x"c9",x"c2"),
  2092 => (x"c9",x"c2",x"78",x"c0"),
  2093 => (x"c0",x"05",x"bf",x"d8"),
  2094 => (x"cf",x"c4",x"87",x"f9"),
  2095 => (x"d6",x"f4",x"49",x"f8"),
  2096 => (x"a8",x"b7",x"c0",x"87"),
  2097 => (x"c4",x"87",x"cd",x"04"),
  2098 => (x"f4",x"49",x"f8",x"cf"),
  2099 => (x"b7",x"c0",x"87",x"c9"),
  2100 => (x"87",x"f3",x"03",x"a8"),
  2101 => (x"bf",x"d8",x"c9",x"c2"),
  2102 => (x"d8",x"c9",x"c2",x"49"),
  2103 => (x"78",x"a1",x"c1",x"48"),
  2104 => (x"81",x"e8",x"c9",x"c2"),
  2105 => (x"c9",x"c2",x"48",x"11"),
  2106 => (x"c9",x"c2",x"58",x"e0"),
  2107 => (x"78",x"c0",x"48",x"e0"),
  2108 => (x"c2",x"87",x"d8",x"c5"),
  2109 => (x"02",x"bf",x"e0",x"c9"),
  2110 => (x"c4",x"87",x"f2",x"c1"),
  2111 => (x"f3",x"49",x"f8",x"cf"),
  2112 => (x"b7",x"c0",x"87",x"d5"),
  2113 => (x"87",x"cd",x"04",x"a8"),
  2114 => (x"bf",x"e0",x"c9",x"c2"),
  2115 => (x"c2",x"88",x"c1",x"48"),
  2116 => (x"db",x"58",x"e4",x"c9"),
  2117 => (x"cc",x"d0",x"c4",x"87"),
  2118 => (x"f6",x"c1",x"49",x"bf"),
  2119 => (x"98",x"70",x"87",x"fe"),
  2120 => (x"c4",x"87",x"cd",x"02"),
  2121 => (x"f0",x"49",x"f8",x"cf"),
  2122 => (x"c9",x"c2",x"87",x"e2"),
  2123 => (x"78",x"c0",x"48",x"d8"),
  2124 => (x"bf",x"dc",x"c9",x"c2"),
  2125 => (x"87",x"d3",x"c4",x"05"),
  2126 => (x"bf",x"e0",x"c9",x"c2"),
  2127 => (x"87",x"cb",x"c4",x"05"),
  2128 => (x"bf",x"d8",x"c9",x"c2"),
  2129 => (x"d8",x"c9",x"c2",x"49"),
  2130 => (x"78",x"a1",x"c1",x"48"),
  2131 => (x"81",x"e8",x"c9",x"c2"),
  2132 => (x"c2",x"49",x"4c",x"11"),
  2133 => (x"c0",x"02",x"99",x"c0"),
  2134 => (x"48",x"74",x"87",x"cc"),
  2135 => (x"c2",x"98",x"ff",x"c1"),
  2136 => (x"c3",x"58",x"e4",x"c9"),
  2137 => (x"c9",x"c2",x"87",x"e5"),
  2138 => (x"de",x"c3",x"5c",x"e0"),
  2139 => (x"dc",x"c9",x"c2",x"87"),
  2140 => (x"ff",x"c0",x"02",x"bf"),
  2141 => (x"d8",x"c9",x"c2",x"87"),
  2142 => (x"c9",x"c2",x"49",x"bf"),
  2143 => (x"a1",x"c1",x"48",x"d8"),
  2144 => (x"e8",x"c9",x"c2",x"78"),
  2145 => (x"49",x"69",x"97",x"81"),
  2146 => (x"f8",x"cf",x"c4",x"1e"),
  2147 => (x"87",x"d3",x"ef",x"49"),
  2148 => (x"c9",x"c2",x"86",x"c4"),
  2149 => (x"c1",x"48",x"bf",x"dc"),
  2150 => (x"e0",x"c9",x"c2",x"88"),
  2151 => (x"e0",x"c9",x"c2",x"58"),
  2152 => (x"c0",x"78",x"c1",x"48"),
  2153 => (x"c1",x"49",x"ec",x"f6"),
  2154 => (x"70",x"87",x"e5",x"f4"),
  2155 => (x"d0",x"d0",x"c4",x"49"),
  2156 => (x"87",x"d7",x"c2",x"59"),
  2157 => (x"49",x"f8",x"cf",x"c4"),
  2158 => (x"70",x"87",x"dc",x"f0"),
  2159 => (x"ab",x"b7",x"c0",x"4b"),
  2160 => (x"87",x"c7",x"c2",x"04"),
  2161 => (x"bf",x"d4",x"c9",x"c2"),
  2162 => (x"87",x"e0",x"c0",x"02"),
  2163 => (x"bf",x"cc",x"d0",x"c4"),
  2164 => (x"c7",x"f4",x"c1",x"49"),
  2165 => (x"02",x"98",x"70",x"87"),
  2166 => (x"c7",x"87",x"d1",x"c0"),
  2167 => (x"e4",x"c9",x"c2",x"48"),
  2168 => (x"c9",x"c2",x"88",x"bf"),
  2169 => (x"c9",x"c2",x"58",x"e8"),
  2170 => (x"78",x"c0",x"48",x"d4"),
  2171 => (x"bf",x"d4",x"c9",x"c2"),
  2172 => (x"49",x"a2",x"c1",x"4a"),
  2173 => (x"59",x"d8",x"c9",x"c2"),
  2174 => (x"82",x"d0",x"d0",x"c4"),
  2175 => (x"c9",x"c2",x"52",x"73"),
  2176 => (x"a9",x"b7",x"bf",x"e4"),
  2177 => (x"87",x"e6",x"c0",x"04"),
  2178 => (x"97",x"d0",x"d0",x"c4"),
  2179 => (x"c4",x"1e",x"49",x"bf"),
  2180 => (x"87",x"e4",x"c1",x"49"),
  2181 => (x"d0",x"c4",x"86",x"c4"),
  2182 => (x"7d",x"bf",x"97",x"d1"),
  2183 => (x"97",x"d2",x"d0",x"c4"),
  2184 => (x"d0",x"ff",x"7d",x"bf"),
  2185 => (x"78",x"e0",x"c0",x"48"),
  2186 => (x"48",x"d4",x"c9",x"c2"),
  2187 => (x"f4",x"c7",x"78",x"c0"),
  2188 => (x"db",x"f2",x"c1",x"49"),
  2189 => (x"c4",x"49",x"70",x"87"),
  2190 => (x"c4",x"59",x"d0",x"d0"),
  2191 => (x"ee",x"49",x"f8",x"cf"),
  2192 => (x"4b",x"70",x"87",x"d5"),
  2193 => (x"03",x"ab",x"b7",x"c0"),
  2194 => (x"26",x"87",x"f9",x"fd"),
  2195 => (x"26",x"4c",x"26",x"4d"),
  2196 => (x"00",x"4f",x"26",x"4b"),
  2197 => (x"00",x"00",x"00",x"00"),
  2198 => (x"00",x"00",x"00",x"00"),
  2199 => (x"00",x"00",x"00",x"00"),
  2200 => (x"00",x"00",x"00",x"00"),
  2201 => (x"00",x"00",x"00",x"04"),
  2202 => (x"08",x"82",x"ff",x"01"),
  2203 => (x"64",x"f3",x"c8",x"f3"),
  2204 => (x"01",x"f2",x"50",x"f3"),
  2205 => (x"00",x"f4",x"01",x"81"),
  2206 => (x"48",x"d0",x"ff",x"1e"),
  2207 => (x"71",x"78",x"e1",x"c8"),
  2208 => (x"08",x"d4",x"ff",x"48"),
  2209 => (x"48",x"66",x"c4",x"78"),
  2210 => (x"78",x"08",x"d4",x"ff"),
  2211 => (x"71",x"1e",x"4f",x"26"),
  2212 => (x"49",x"66",x"c4",x"4a"),
  2213 => (x"ff",x"49",x"72",x"1e"),
  2214 => (x"d0",x"ff",x"87",x"de"),
  2215 => (x"78",x"e0",x"c0",x"48"),
  2216 => (x"4f",x"26",x"8e",x"fc"),
  2217 => (x"71",x"1e",x"73",x"1e"),
  2218 => (x"49",x"66",x"c8",x"4b"),
  2219 => (x"c1",x"4a",x"73",x"1e"),
  2220 => (x"ff",x"49",x"a2",x"e0"),
  2221 => (x"8e",x"fc",x"87",x"d8"),
  2222 => (x"4f",x"26",x"4b",x"26"),
  2223 => (x"4a",x"d4",x"ff",x"1e"),
  2224 => (x"ff",x"7a",x"ff",x"c3"),
  2225 => (x"e1",x"c0",x"48",x"d0"),
  2226 => (x"c4",x"7a",x"de",x"78"),
  2227 => (x"7a",x"bf",x"d4",x"d0"),
  2228 => (x"28",x"c8",x"48",x"49"),
  2229 => (x"48",x"71",x"7a",x"70"),
  2230 => (x"7a",x"70",x"28",x"d0"),
  2231 => (x"28",x"d8",x"48",x"71"),
  2232 => (x"d0",x"ff",x"7a",x"70"),
  2233 => (x"78",x"e0",x"c0",x"48"),
  2234 => (x"5e",x"0e",x"4f",x"26"),
  2235 => (x"0e",x"5d",x"5c",x"5b"),
  2236 => (x"d0",x"c4",x"4c",x"71"),
  2237 => (x"49",x"4d",x"bf",x"d4"),
  2238 => (x"4b",x"71",x"29",x"74"),
  2239 => (x"c1",x"9b",x"66",x"d0"),
  2240 => (x"b7",x"66",x"d4",x"83"),
  2241 => (x"87",x"c2",x"04",x"ab"),
  2242 => (x"66",x"d0",x"4b",x"c0"),
  2243 => (x"ff",x"31",x"74",x"49"),
  2244 => (x"73",x"99",x"75",x"b9"),
  2245 => (x"72",x"32",x"74",x"4a"),
  2246 => (x"c4",x"b0",x"71",x"48"),
  2247 => (x"fe",x"58",x"d8",x"d0"),
  2248 => (x"4d",x"26",x"87",x"da"),
  2249 => (x"4b",x"26",x"4c",x"26"),
  2250 => (x"ff",x"1e",x"4f",x"26"),
  2251 => (x"c9",x"c8",x"48",x"d0"),
  2252 => (x"ff",x"48",x"71",x"78"),
  2253 => (x"26",x"78",x"08",x"d4"),
  2254 => (x"4a",x"71",x"1e",x"4f"),
  2255 => (x"ff",x"87",x"eb",x"49"),
  2256 => (x"78",x"c8",x"48",x"d0"),
  2257 => (x"73",x"1e",x"4f",x"26"),
  2258 => (x"c4",x"4b",x"71",x"1e"),
  2259 => (x"02",x"bf",x"e4",x"d0"),
  2260 => (x"eb",x"c2",x"87",x"c3"),
  2261 => (x"48",x"d0",x"ff",x"87"),
  2262 => (x"73",x"78",x"c9",x"c8"),
  2263 => (x"b1",x"e0",x"c0",x"49"),
  2264 => (x"71",x"48",x"d4",x"ff"),
  2265 => (x"d8",x"d0",x"c4",x"78"),
  2266 => (x"c8",x"78",x"c0",x"48"),
  2267 => (x"87",x"c5",x"02",x"66"),
  2268 => (x"c2",x"49",x"ff",x"c3"),
  2269 => (x"c4",x"49",x"c0",x"87"),
  2270 => (x"cc",x"59",x"e0",x"d0"),
  2271 => (x"87",x"c6",x"02",x"66"),
  2272 => (x"4a",x"d5",x"d5",x"c5"),
  2273 => (x"ff",x"cf",x"87",x"c4"),
  2274 => (x"d0",x"c4",x"4a",x"ff"),
  2275 => (x"d0",x"c4",x"5a",x"e4"),
  2276 => (x"78",x"c1",x"48",x"e4"),
  2277 => (x"4f",x"26",x"4b",x"26"),
  2278 => (x"5c",x"5b",x"5e",x"0e"),
  2279 => (x"4d",x"71",x"0e",x"5d"),
  2280 => (x"bf",x"e0",x"d0",x"c4"),
  2281 => (x"02",x"9d",x"75",x"4b"),
  2282 => (x"c8",x"49",x"87",x"cb"),
  2283 => (x"fc",x"cc",x"c2",x"91"),
  2284 => (x"c4",x"82",x"71",x"4a"),
  2285 => (x"fc",x"d0",x"c2",x"87"),
  2286 => (x"12",x"4c",x"c0",x"4a"),
  2287 => (x"c4",x"99",x"73",x"49"),
  2288 => (x"b9",x"bf",x"dc",x"d0"),
  2289 => (x"71",x"48",x"d4",x"ff"),
  2290 => (x"2b",x"b7",x"c1",x"78"),
  2291 => (x"ac",x"b7",x"c8",x"84"),
  2292 => (x"c4",x"87",x"e8",x"04"),
  2293 => (x"48",x"bf",x"d8",x"d0"),
  2294 => (x"d0",x"c4",x"80",x"c8"),
  2295 => (x"4d",x"26",x"58",x"dc"),
  2296 => (x"4b",x"26",x"4c",x"26"),
  2297 => (x"73",x"1e",x"4f",x"26"),
  2298 => (x"13",x"4b",x"71",x"1e"),
  2299 => (x"cb",x"02",x"9a",x"4a"),
  2300 => (x"fe",x"49",x"72",x"87"),
  2301 => (x"4a",x"13",x"87",x"e2"),
  2302 => (x"87",x"f5",x"05",x"9a"),
  2303 => (x"4f",x"26",x"4b",x"26"),
  2304 => (x"d8",x"d0",x"c4",x"1e"),
  2305 => (x"d0",x"c4",x"49",x"bf"),
  2306 => (x"a1",x"c1",x"48",x"d8"),
  2307 => (x"b7",x"c0",x"c4",x"78"),
  2308 => (x"87",x"db",x"03",x"a9"),
  2309 => (x"c4",x"48",x"d4",x"ff"),
  2310 => (x"78",x"bf",x"dc",x"d0"),
  2311 => (x"bf",x"d8",x"d0",x"c4"),
  2312 => (x"d8",x"d0",x"c4",x"49"),
  2313 => (x"78",x"a1",x"c1",x"48"),
  2314 => (x"a9",x"b7",x"c0",x"c4"),
  2315 => (x"ff",x"87",x"e5",x"04"),
  2316 => (x"78",x"c8",x"48",x"d0"),
  2317 => (x"48",x"e4",x"d0",x"c4"),
  2318 => (x"4f",x"26",x"78",x"c0"),
  2319 => (x"00",x"00",x"00",x"00"),
  2320 => (x"00",x"00",x"00",x"00"),
  2321 => (x"5f",x"00",x"00",x"00"),
  2322 => (x"00",x"00",x"00",x"5f"),
  2323 => (x"00",x"03",x"03",x"00"),
  2324 => (x"00",x"00",x"03",x"03"),
  2325 => (x"14",x"7f",x"7f",x"14"),
  2326 => (x"00",x"14",x"7f",x"7f"),
  2327 => (x"6b",x"2e",x"24",x"00"),
  2328 => (x"00",x"12",x"3a",x"6b"),
  2329 => (x"18",x"36",x"6a",x"4c"),
  2330 => (x"00",x"32",x"56",x"6c"),
  2331 => (x"59",x"4f",x"7e",x"30"),
  2332 => (x"40",x"68",x"3a",x"77"),
  2333 => (x"07",x"04",x"00",x"00"),
  2334 => (x"00",x"00",x"00",x"03"),
  2335 => (x"3e",x"1c",x"00",x"00"),
  2336 => (x"00",x"00",x"41",x"63"),
  2337 => (x"63",x"41",x"00",x"00"),
  2338 => (x"00",x"00",x"1c",x"3e"),
  2339 => (x"1c",x"3e",x"2a",x"08"),
  2340 => (x"08",x"2a",x"3e",x"1c"),
  2341 => (x"3e",x"08",x"08",x"00"),
  2342 => (x"00",x"08",x"08",x"3e"),
  2343 => (x"e0",x"80",x"00",x"00"),
  2344 => (x"00",x"00",x"00",x"60"),
  2345 => (x"08",x"08",x"08",x"00"),
  2346 => (x"00",x"08",x"08",x"08"),
  2347 => (x"60",x"00",x"00",x"00"),
  2348 => (x"00",x"00",x"00",x"60"),
  2349 => (x"18",x"30",x"60",x"40"),
  2350 => (x"01",x"03",x"06",x"0c"),
  2351 => (x"59",x"7f",x"3e",x"00"),
  2352 => (x"00",x"3e",x"7f",x"4d"),
  2353 => (x"7f",x"06",x"04",x"00"),
  2354 => (x"00",x"00",x"00",x"7f"),
  2355 => (x"71",x"63",x"42",x"00"),
  2356 => (x"00",x"46",x"4f",x"59"),
  2357 => (x"49",x"63",x"22",x"00"),
  2358 => (x"00",x"36",x"7f",x"49"),
  2359 => (x"13",x"16",x"1c",x"18"),
  2360 => (x"00",x"10",x"7f",x"7f"),
  2361 => (x"45",x"67",x"27",x"00"),
  2362 => (x"00",x"39",x"7d",x"45"),
  2363 => (x"4b",x"7e",x"3c",x"00"),
  2364 => (x"00",x"30",x"79",x"49"),
  2365 => (x"71",x"01",x"01",x"00"),
  2366 => (x"00",x"07",x"0f",x"79"),
  2367 => (x"49",x"7f",x"36",x"00"),
  2368 => (x"00",x"36",x"7f",x"49"),
  2369 => (x"49",x"4f",x"06",x"00"),
  2370 => (x"00",x"1e",x"3f",x"69"),
  2371 => (x"66",x"00",x"00",x"00"),
  2372 => (x"00",x"00",x"00",x"66"),
  2373 => (x"e6",x"80",x"00",x"00"),
  2374 => (x"00",x"00",x"00",x"66"),
  2375 => (x"14",x"08",x"08",x"00"),
  2376 => (x"00",x"22",x"22",x"14"),
  2377 => (x"14",x"14",x"14",x"00"),
  2378 => (x"00",x"14",x"14",x"14"),
  2379 => (x"14",x"22",x"22",x"00"),
  2380 => (x"00",x"08",x"08",x"14"),
  2381 => (x"51",x"03",x"02",x"00"),
  2382 => (x"00",x"06",x"0f",x"59"),
  2383 => (x"5d",x"41",x"7f",x"3e"),
  2384 => (x"00",x"1e",x"1f",x"55"),
  2385 => (x"09",x"7f",x"7e",x"00"),
  2386 => (x"00",x"7e",x"7f",x"09"),
  2387 => (x"49",x"7f",x"7f",x"00"),
  2388 => (x"00",x"36",x"7f",x"49"),
  2389 => (x"63",x"3e",x"1c",x"00"),
  2390 => (x"00",x"41",x"41",x"41"),
  2391 => (x"41",x"7f",x"7f",x"00"),
  2392 => (x"00",x"1c",x"3e",x"63"),
  2393 => (x"49",x"7f",x"7f",x"00"),
  2394 => (x"00",x"41",x"41",x"49"),
  2395 => (x"09",x"7f",x"7f",x"00"),
  2396 => (x"00",x"01",x"01",x"09"),
  2397 => (x"41",x"7f",x"3e",x"00"),
  2398 => (x"00",x"7a",x"7b",x"49"),
  2399 => (x"08",x"7f",x"7f",x"00"),
  2400 => (x"00",x"7f",x"7f",x"08"),
  2401 => (x"7f",x"41",x"00",x"00"),
  2402 => (x"00",x"00",x"41",x"7f"),
  2403 => (x"40",x"60",x"20",x"00"),
  2404 => (x"00",x"3f",x"7f",x"40"),
  2405 => (x"1c",x"08",x"7f",x"7f"),
  2406 => (x"00",x"41",x"63",x"36"),
  2407 => (x"40",x"7f",x"7f",x"00"),
  2408 => (x"00",x"40",x"40",x"40"),
  2409 => (x"0c",x"06",x"7f",x"7f"),
  2410 => (x"00",x"7f",x"7f",x"06"),
  2411 => (x"0c",x"06",x"7f",x"7f"),
  2412 => (x"00",x"7f",x"7f",x"18"),
  2413 => (x"41",x"7f",x"3e",x"00"),
  2414 => (x"00",x"3e",x"7f",x"41"),
  2415 => (x"09",x"7f",x"7f",x"00"),
  2416 => (x"00",x"06",x"0f",x"09"),
  2417 => (x"61",x"41",x"7f",x"3e"),
  2418 => (x"00",x"40",x"7e",x"7f"),
  2419 => (x"09",x"7f",x"7f",x"00"),
  2420 => (x"00",x"66",x"7f",x"19"),
  2421 => (x"4d",x"6f",x"26",x"00"),
  2422 => (x"00",x"32",x"7b",x"59"),
  2423 => (x"7f",x"01",x"01",x"00"),
  2424 => (x"00",x"01",x"01",x"7f"),
  2425 => (x"40",x"7f",x"3f",x"00"),
  2426 => (x"00",x"3f",x"7f",x"40"),
  2427 => (x"70",x"3f",x"0f",x"00"),
  2428 => (x"00",x"0f",x"3f",x"70"),
  2429 => (x"18",x"30",x"7f",x"7f"),
  2430 => (x"00",x"7f",x"7f",x"30"),
  2431 => (x"1c",x"36",x"63",x"41"),
  2432 => (x"41",x"63",x"36",x"1c"),
  2433 => (x"7c",x"06",x"03",x"01"),
  2434 => (x"01",x"03",x"06",x"7c"),
  2435 => (x"4d",x"59",x"71",x"61"),
  2436 => (x"00",x"41",x"43",x"47"),
  2437 => (x"7f",x"7f",x"00",x"00"),
  2438 => (x"00",x"00",x"41",x"41"),
  2439 => (x"0c",x"06",x"03",x"01"),
  2440 => (x"40",x"60",x"30",x"18"),
  2441 => (x"41",x"41",x"00",x"00"),
  2442 => (x"00",x"00",x"7f",x"7f"),
  2443 => (x"03",x"06",x"0c",x"08"),
  2444 => (x"00",x"08",x"0c",x"06"),
  2445 => (x"80",x"80",x"80",x"80"),
  2446 => (x"00",x"80",x"80",x"80"),
  2447 => (x"03",x"00",x"00",x"00"),
  2448 => (x"00",x"00",x"04",x"07"),
  2449 => (x"54",x"74",x"20",x"00"),
  2450 => (x"00",x"78",x"7c",x"54"),
  2451 => (x"44",x"7f",x"7f",x"00"),
  2452 => (x"00",x"38",x"7c",x"44"),
  2453 => (x"44",x"7c",x"38",x"00"),
  2454 => (x"00",x"00",x"44",x"44"),
  2455 => (x"44",x"7c",x"38",x"00"),
  2456 => (x"00",x"7f",x"7f",x"44"),
  2457 => (x"54",x"7c",x"38",x"00"),
  2458 => (x"00",x"18",x"5c",x"54"),
  2459 => (x"7f",x"7e",x"04",x"00"),
  2460 => (x"00",x"00",x"05",x"05"),
  2461 => (x"a4",x"bc",x"18",x"00"),
  2462 => (x"00",x"7c",x"fc",x"a4"),
  2463 => (x"04",x"7f",x"7f",x"00"),
  2464 => (x"00",x"78",x"7c",x"04"),
  2465 => (x"3d",x"00",x"00",x"00"),
  2466 => (x"00",x"00",x"40",x"7d"),
  2467 => (x"80",x"80",x"80",x"00"),
  2468 => (x"00",x"00",x"7d",x"fd"),
  2469 => (x"10",x"7f",x"7f",x"00"),
  2470 => (x"00",x"44",x"6c",x"38"),
  2471 => (x"3f",x"00",x"00",x"00"),
  2472 => (x"00",x"00",x"40",x"7f"),
  2473 => (x"18",x"0c",x"7c",x"7c"),
  2474 => (x"00",x"78",x"7c",x"0c"),
  2475 => (x"04",x"7c",x"7c",x"00"),
  2476 => (x"00",x"78",x"7c",x"04"),
  2477 => (x"44",x"7c",x"38",x"00"),
  2478 => (x"00",x"38",x"7c",x"44"),
  2479 => (x"24",x"fc",x"fc",x"00"),
  2480 => (x"00",x"18",x"3c",x"24"),
  2481 => (x"24",x"3c",x"18",x"00"),
  2482 => (x"00",x"fc",x"fc",x"24"),
  2483 => (x"04",x"7c",x"7c",x"00"),
  2484 => (x"00",x"08",x"0c",x"04"),
  2485 => (x"54",x"5c",x"48",x"00"),
  2486 => (x"00",x"20",x"74",x"54"),
  2487 => (x"7f",x"3f",x"04",x"00"),
  2488 => (x"00",x"00",x"44",x"44"),
  2489 => (x"40",x"7c",x"3c",x"00"),
  2490 => (x"00",x"7c",x"7c",x"40"),
  2491 => (x"60",x"3c",x"1c",x"00"),
  2492 => (x"00",x"1c",x"3c",x"60"),
  2493 => (x"30",x"60",x"7c",x"3c"),
  2494 => (x"00",x"3c",x"7c",x"60"),
  2495 => (x"10",x"38",x"6c",x"44"),
  2496 => (x"00",x"44",x"6c",x"38"),
  2497 => (x"e0",x"bc",x"1c",x"00"),
  2498 => (x"00",x"1c",x"3c",x"60"),
  2499 => (x"74",x"64",x"44",x"00"),
  2500 => (x"00",x"44",x"4c",x"5c"),
  2501 => (x"3e",x"08",x"08",x"00"),
  2502 => (x"00",x"41",x"41",x"77"),
  2503 => (x"7f",x"00",x"00",x"00"),
  2504 => (x"00",x"00",x"00",x"7f"),
  2505 => (x"77",x"41",x"41",x"00"),
  2506 => (x"00",x"08",x"08",x"3e"),
  2507 => (x"03",x"01",x"01",x"02"),
  2508 => (x"00",x"01",x"02",x"02"),
  2509 => (x"7f",x"7f",x"7f",x"7f"),
  2510 => (x"00",x"7f",x"7f",x"7f"),
  2511 => (x"1c",x"1c",x"08",x"08"),
  2512 => (x"7f",x"7f",x"3e",x"3e"),
  2513 => (x"3e",x"3e",x"7f",x"7f"),
  2514 => (x"08",x"08",x"1c",x"1c"),
  2515 => (x"7c",x"18",x"10",x"00"),
  2516 => (x"00",x"10",x"18",x"7c"),
  2517 => (x"7c",x"30",x"10",x"00"),
  2518 => (x"00",x"10",x"30",x"7c"),
  2519 => (x"60",x"60",x"30",x"10"),
  2520 => (x"00",x"06",x"1e",x"78"),
  2521 => (x"18",x"3c",x"66",x"42"),
  2522 => (x"00",x"42",x"66",x"3c"),
  2523 => (x"c2",x"6a",x"38",x"78"),
  2524 => (x"00",x"38",x"6c",x"c6"),
  2525 => (x"60",x"00",x"00",x"60"),
  2526 => (x"00",x"60",x"00",x"00"),
  2527 => (x"5c",x"5b",x"5e",x"0e"),
  2528 => (x"86",x"fc",x"0e",x"5d"),
  2529 => (x"d0",x"c4",x"7e",x"71"),
  2530 => (x"c0",x"4c",x"bf",x"f8"),
  2531 => (x"c4",x"1e",x"c0",x"4b"),
  2532 => (x"c4",x"02",x"ab",x"66"),
  2533 => (x"c2",x"4d",x"c0",x"87"),
  2534 => (x"75",x"4d",x"c1",x"87"),
  2535 => (x"ee",x"49",x"73",x"1e"),
  2536 => (x"86",x"c8",x"87",x"e4"),
  2537 => (x"ef",x"49",x"e0",x"c0"),
  2538 => (x"a4",x"c4",x"87",x"ee"),
  2539 => (x"f0",x"49",x"6a",x"4a"),
  2540 => (x"cb",x"f1",x"87",x"f4"),
  2541 => (x"c1",x"84",x"cc",x"87"),
  2542 => (x"ab",x"b7",x"c8",x"83"),
  2543 => (x"87",x"cd",x"ff",x"04"),
  2544 => (x"4d",x"26",x"8e",x"fc"),
  2545 => (x"4b",x"26",x"4c",x"26"),
  2546 => (x"71",x"1e",x"4f",x"26"),
  2547 => (x"fc",x"d0",x"c4",x"4a"),
  2548 => (x"fc",x"d0",x"c4",x"5a"),
  2549 => (x"49",x"78",x"c7",x"48"),
  2550 => (x"26",x"87",x"e1",x"fe"),
  2551 => (x"1e",x"73",x"1e",x"4f"),
  2552 => (x"b7",x"c0",x"4a",x"71"),
  2553 => (x"87",x"d3",x"03",x"aa"),
  2554 => (x"bf",x"e0",x"ee",x"c2"),
  2555 => (x"c1",x"87",x"c4",x"05"),
  2556 => (x"c0",x"87",x"c2",x"4b"),
  2557 => (x"e4",x"ee",x"c2",x"4b"),
  2558 => (x"c2",x"87",x"c4",x"5b"),
  2559 => (x"c2",x"5a",x"e4",x"ee"),
  2560 => (x"4a",x"bf",x"e0",x"ee"),
  2561 => (x"c0",x"c1",x"9a",x"c1"),
  2562 => (x"ec",x"ec",x"49",x"a2"),
  2563 => (x"c2",x"48",x"fc",x"87"),
  2564 => (x"78",x"bf",x"e0",x"ee"),
  2565 => (x"4f",x"26",x"4b",x"26"),
  2566 => (x"c4",x"4a",x"71",x"1e"),
  2567 => (x"49",x"72",x"1e",x"66"),
  2568 => (x"fc",x"87",x"c1",x"ea"),
  2569 => (x"1e",x"4f",x"26",x"8e"),
  2570 => (x"bf",x"e0",x"ee",x"c2"),
  2571 => (x"cb",x"df",x"ff",x"49"),
  2572 => (x"f0",x"d0",x"c4",x"87"),
  2573 => (x"78",x"bf",x"e8",x"48"),
  2574 => (x"48",x"ec",x"d0",x"c4"),
  2575 => (x"c4",x"78",x"bf",x"ec"),
  2576 => (x"4a",x"bf",x"f0",x"d0"),
  2577 => (x"99",x"ff",x"c3",x"49"),
  2578 => (x"72",x"2a",x"b7",x"c8"),
  2579 => (x"c4",x"b0",x"71",x"48"),
  2580 => (x"26",x"58",x"f8",x"d0"),
  2581 => (x"5b",x"5e",x"0e",x"4f"),
  2582 => (x"71",x"0e",x"5d",x"5c"),
  2583 => (x"87",x"c7",x"ff",x"4b"),
  2584 => (x"48",x"e8",x"d0",x"c4"),
  2585 => (x"49",x"73",x"50",x"c0"),
  2586 => (x"87",x"f0",x"de",x"ff"),
  2587 => (x"c2",x"4c",x"49",x"70"),
  2588 => (x"49",x"ee",x"cb",x"9c"),
  2589 => (x"87",x"d8",x"d9",x"c1"),
  2590 => (x"c4",x"4d",x"49",x"70"),
  2591 => (x"bf",x"97",x"e8",x"d0"),
  2592 => (x"87",x"e5",x"c1",x"05"),
  2593 => (x"c4",x"49",x"66",x"d0"),
  2594 => (x"99",x"bf",x"f4",x"d0"),
  2595 => (x"d4",x"87",x"d7",x"05"),
  2596 => (x"d0",x"c4",x"49",x"66"),
  2597 => (x"05",x"99",x"bf",x"ec"),
  2598 => (x"49",x"73",x"87",x"cc"),
  2599 => (x"87",x"fc",x"dd",x"ff"),
  2600 => (x"c1",x"02",x"98",x"70"),
  2601 => (x"4c",x"c1",x"87",x"c3"),
  2602 => (x"75",x"87",x"fc",x"fd"),
  2603 => (x"eb",x"d8",x"c1",x"49"),
  2604 => (x"02",x"98",x"70",x"87"),
  2605 => (x"d0",x"c4",x"87",x"c6"),
  2606 => (x"50",x"c1",x"48",x"e8"),
  2607 => (x"97",x"e8",x"d0",x"c4"),
  2608 => (x"e4",x"c0",x"05",x"bf"),
  2609 => (x"f4",x"d0",x"c4",x"87"),
  2610 => (x"66",x"d0",x"49",x"bf"),
  2611 => (x"d5",x"ff",x"05",x"99"),
  2612 => (x"ec",x"d0",x"c4",x"87"),
  2613 => (x"66",x"d4",x"49",x"bf"),
  2614 => (x"c9",x"ff",x"05",x"99"),
  2615 => (x"ff",x"49",x"73",x"87"),
  2616 => (x"70",x"87",x"f9",x"dc"),
  2617 => (x"fd",x"fe",x"05",x"98"),
  2618 => (x"26",x"48",x"74",x"87"),
  2619 => (x"26",x"4c",x"26",x"4d"),
  2620 => (x"0e",x"4f",x"26",x"4b"),
  2621 => (x"5d",x"5c",x"5b",x"5e"),
  2622 => (x"c8",x"86",x"f0",x"0e"),
  2623 => (x"78",x"c0",x"48",x"a6"),
  2624 => (x"78",x"c0",x"80",x"c4"),
  2625 => (x"f8",x"7e",x"bf",x"ec"),
  2626 => (x"f8",x"d0",x"c4",x"80"),
  2627 => (x"1e",x"c1",x"78",x"bf"),
  2628 => (x"49",x"c7",x"1e",x"c0"),
  2629 => (x"c8",x"87",x"fe",x"fc"),
  2630 => (x"02",x"98",x"70",x"86"),
  2631 => (x"49",x"ff",x"87",x"d1"),
  2632 => (x"c1",x"87",x"fa",x"fa"),
  2633 => (x"db",x"ff",x"49",x"da"),
  2634 => (x"a6",x"c8",x"87",x"f2"),
  2635 => (x"c4",x"78",x"c1",x"48"),
  2636 => (x"bf",x"97",x"e8",x"d0"),
  2637 => (x"c1",x"87",x"c4",x"02"),
  2638 => (x"c4",x"87",x"fa",x"d6"),
  2639 => (x"4b",x"bf",x"f0",x"d0"),
  2640 => (x"bf",x"e0",x"ee",x"c2"),
  2641 => (x"87",x"c7",x"c1",x"05"),
  2642 => (x"4d",x"c0",x"c0",x"c8"),
  2643 => (x"4c",x"e4",x"fd",x"c3"),
  2644 => (x"db",x"ff",x"49",x"14"),
  2645 => (x"98",x"70",x"87",x"c6"),
  2646 => (x"75",x"87",x"c2",x"02"),
  2647 => (x"2d",x"b7",x"c1",x"b3"),
  2648 => (x"87",x"ec",x"ff",x"05"),
  2649 => (x"ff",x"49",x"fd",x"c3"),
  2650 => (x"c3",x"87",x"f1",x"da"),
  2651 => (x"da",x"ff",x"49",x"fa"),
  2652 => (x"49",x"73",x"87",x"ea"),
  2653 => (x"71",x"99",x"ff",x"c3"),
  2654 => (x"fa",x"49",x"c0",x"1e"),
  2655 => (x"49",x"73",x"87",x"da"),
  2656 => (x"71",x"29",x"b7",x"c8"),
  2657 => (x"fa",x"49",x"c1",x"1e"),
  2658 => (x"86",x"c8",x"87",x"ce"),
  2659 => (x"c4",x"87",x"e9",x"c6"),
  2660 => (x"4b",x"bf",x"f4",x"d0"),
  2661 => (x"e0",x"c0",x"02",x"9b"),
  2662 => (x"dc",x"ee",x"c2",x"87"),
  2663 => (x"d4",x"c1",x"49",x"bf"),
  2664 => (x"98",x"70",x"87",x"fa"),
  2665 => (x"c0",x"87",x"c4",x"05"),
  2666 => (x"c2",x"87",x"d4",x"4b"),
  2667 => (x"d4",x"c1",x"49",x"e0"),
  2668 => (x"ee",x"c2",x"87",x"de"),
  2669 => (x"c6",x"c0",x"58",x"e0"),
  2670 => (x"dc",x"ee",x"c2",x"87"),
  2671 => (x"73",x"78",x"c0",x"48"),
  2672 => (x"05",x"99",x"c2",x"49"),
  2673 => (x"eb",x"c3",x"87",x"cf"),
  2674 => (x"cf",x"d9",x"ff",x"49"),
  2675 => (x"c2",x"49",x"70",x"87"),
  2676 => (x"c5",x"c0",x"02",x"99"),
  2677 => (x"48",x"a6",x"cc",x"87"),
  2678 => (x"49",x"73",x"78",x"fb"),
  2679 => (x"cf",x"05",x"99",x"c1"),
  2680 => (x"49",x"f4",x"c3",x"87"),
  2681 => (x"87",x"f4",x"d8",x"ff"),
  2682 => (x"99",x"c2",x"49",x"70"),
  2683 => (x"87",x"c5",x"c0",x"02"),
  2684 => (x"fa",x"48",x"a6",x"cc"),
  2685 => (x"c8",x"49",x"73",x"78"),
  2686 => (x"ce",x"c0",x"05",x"99"),
  2687 => (x"49",x"f5",x"c3",x"87"),
  2688 => (x"87",x"d8",x"d8",x"ff"),
  2689 => (x"99",x"c2",x"49",x"70"),
  2690 => (x"c4",x"87",x"dc",x"02"),
  2691 => (x"02",x"bf",x"fc",x"d0"),
  2692 => (x"48",x"87",x"ca",x"c0"),
  2693 => (x"d1",x"c4",x"88",x"c1"),
  2694 => (x"c5",x"c0",x"58",x"c0"),
  2695 => (x"48",x"a6",x"cc",x"87"),
  2696 => (x"a6",x"c8",x"78",x"ff"),
  2697 => (x"73",x"78",x"c1",x"48"),
  2698 => (x"05",x"99",x"c4",x"49"),
  2699 => (x"c3",x"87",x"cf",x"c0"),
  2700 => (x"d7",x"ff",x"49",x"f2"),
  2701 => (x"49",x"70",x"87",x"e6"),
  2702 => (x"c0",x"02",x"99",x"c2"),
  2703 => (x"d0",x"c4",x"87",x"e2"),
  2704 => (x"48",x"7e",x"bf",x"fc"),
  2705 => (x"03",x"a8",x"b7",x"c7"),
  2706 => (x"6e",x"87",x"cb",x"c0"),
  2707 => (x"c4",x"80",x"c1",x"48"),
  2708 => (x"c0",x"58",x"c0",x"d1"),
  2709 => (x"a6",x"cc",x"87",x"c5"),
  2710 => (x"c8",x"78",x"fe",x"48"),
  2711 => (x"78",x"c1",x"48",x"a6"),
  2712 => (x"ff",x"49",x"fd",x"c3"),
  2713 => (x"70",x"87",x"f5",x"d6"),
  2714 => (x"02",x"99",x"c2",x"49"),
  2715 => (x"c4",x"87",x"db",x"c0"),
  2716 => (x"02",x"bf",x"fc",x"d0"),
  2717 => (x"c4",x"87",x"c9",x"c0"),
  2718 => (x"c0",x"48",x"fc",x"d0"),
  2719 => (x"87",x"c5",x"c0",x"78"),
  2720 => (x"fd",x"48",x"a6",x"cc"),
  2721 => (x"48",x"a6",x"c8",x"78"),
  2722 => (x"fa",x"c3",x"78",x"c1"),
  2723 => (x"cb",x"d6",x"ff",x"49"),
  2724 => (x"c2",x"49",x"70",x"87"),
  2725 => (x"df",x"c0",x"02",x"99"),
  2726 => (x"fc",x"d0",x"c4",x"87"),
  2727 => (x"b7",x"c7",x"48",x"bf"),
  2728 => (x"c9",x"c0",x"03",x"a8"),
  2729 => (x"fc",x"d0",x"c4",x"87"),
  2730 => (x"c0",x"78",x"c7",x"48"),
  2731 => (x"a6",x"cc",x"87",x"c5"),
  2732 => (x"c8",x"78",x"fc",x"48"),
  2733 => (x"78",x"c1",x"48",x"a6"),
  2734 => (x"c0",x"48",x"66",x"cc"),
  2735 => (x"c0",x"03",x"a8",x"b7"),
  2736 => (x"66",x"c4",x"87",x"d6"),
  2737 => (x"80",x"e0",x"c1",x"48"),
  2738 => (x"bf",x"6e",x"7e",x"70"),
  2739 => (x"87",x"c8",x"c0",x"02"),
  2740 => (x"cc",x"4b",x"bf",x"6e"),
  2741 => (x"0f",x"73",x"49",x"66"),
  2742 => (x"f0",x"c3",x"1e",x"c0"),
  2743 => (x"49",x"da",x"c1",x"1e"),
  2744 => (x"c8",x"87",x"f2",x"f5"),
  2745 => (x"02",x"98",x"70",x"86"),
  2746 => (x"c4",x"87",x"d9",x"c0"),
  2747 => (x"7e",x"bf",x"fc",x"d0"),
  2748 => (x"91",x"cc",x"49",x"6e"),
  2749 => (x"71",x"4a",x"66",x"c4"),
  2750 => (x"c0",x"02",x"6a",x"82"),
  2751 => (x"4b",x"6a",x"87",x"c6"),
  2752 => (x"0f",x"73",x"49",x"6e"),
  2753 => (x"c0",x"02",x"66",x"c8"),
  2754 => (x"d0",x"c4",x"87",x"c8"),
  2755 => (x"f1",x"49",x"bf",x"fc"),
  2756 => (x"ee",x"c2",x"87",x"ea"),
  2757 => (x"c0",x"02",x"bf",x"e4"),
  2758 => (x"c1",x"49",x"87",x"de"),
  2759 => (x"70",x"87",x"fd",x"ce"),
  2760 => (x"d3",x"c0",x"02",x"98"),
  2761 => (x"fc",x"d0",x"c4",x"87"),
  2762 => (x"cf",x"f1",x"49",x"bf"),
  2763 => (x"f2",x"49",x"c0",x"87"),
  2764 => (x"ee",x"c2",x"87",x"eb"),
  2765 => (x"78",x"c0",x"48",x"e4"),
  2766 => (x"4d",x"26",x"8e",x"f0"),
  2767 => (x"4b",x"26",x"4c",x"26"),
  2768 => (x"5e",x"0e",x"4f",x"26"),
  2769 => (x"0e",x"5d",x"5c",x"5b"),
  2770 => (x"4c",x"71",x"86",x"fc"),
  2771 => (x"bf",x"f8",x"d0",x"c4"),
  2772 => (x"a1",x"d4",x"c1",x"49"),
  2773 => (x"81",x"d8",x"c1",x"4d"),
  2774 => (x"9c",x"74",x"7e",x"69"),
  2775 => (x"c4",x"87",x"cf",x"02"),
  2776 => (x"7b",x"74",x"4b",x"a5"),
  2777 => (x"bf",x"f8",x"d0",x"c4"),
  2778 => (x"87",x"de",x"f1",x"49"),
  2779 => (x"9c",x"74",x"7b",x"6e"),
  2780 => (x"c0",x"87",x"c4",x"05"),
  2781 => (x"c1",x"87",x"c2",x"4b"),
  2782 => (x"f1",x"49",x"73",x"4b"),
  2783 => (x"66",x"d4",x"87",x"df"),
  2784 => (x"49",x"87",x"c9",x"02"),
  2785 => (x"87",x"c8",x"cd",x"c1"),
  2786 => (x"87",x"c2",x"4a",x"70"),
  2787 => (x"ee",x"c2",x"4a",x"c0"),
  2788 => (x"8e",x"fc",x"5a",x"e8"),
  2789 => (x"4c",x"26",x"4d",x"26"),
  2790 => (x"4f",x"26",x"4b",x"26"),
  2791 => (x"00",x"00",x"00",x"00"),
  2792 => (x"00",x"00",x"00",x"00"),
  2793 => (x"00",x"00",x"00",x"00"),
  2794 => (x"71",x"1e",x"73",x"1e"),
  2795 => (x"cb",x"c1",x"49",x"4b"),
  2796 => (x"d1",x"da",x"fd",x"4a"),
  2797 => (x"1e",x"4a",x"70",x"87"),
  2798 => (x"fc",x"c0",x"49",x"72"),
  2799 => (x"c5",x"da",x"fd",x"4a"),
  2800 => (x"26",x"49",x"70",x"87"),
  2801 => (x"48",x"66",x"c8",x"4a"),
  2802 => (x"49",x"72",x"50",x"71"),
  2803 => (x"fd",x"4a",x"fc",x"c0"),
  2804 => (x"71",x"87",x"f3",x"d9"),
  2805 => (x"49",x"66",x"c8",x"4a"),
  2806 => (x"51",x"72",x"81",x"c1"),
  2807 => (x"cb",x"c1",x"49",x"73"),
  2808 => (x"e1",x"d9",x"fd",x"4a"),
  2809 => (x"c8",x"4a",x"71",x"87"),
  2810 => (x"81",x"c2",x"49",x"66"),
  2811 => (x"4b",x"26",x"51",x"72"),
  2812 => (x"73",x"1e",x"4f",x"26"),
  2813 => (x"c8",x"4b",x"71",x"1e"),
  2814 => (x"cb",x"c1",x"49",x"66"),
  2815 => (x"4a",x"66",x"cc",x"91"),
  2816 => (x"4a",x"73",x"49",x"a1"),
  2817 => (x"92",x"d4",x"c6",x"c1"),
  2818 => (x"c2",x"49",x"a1",x"72"),
  2819 => (x"48",x"71",x"89",x"d6"),
  2820 => (x"4f",x"26",x"4b",x"26"),
  2821 => (x"5c",x"5b",x"5e",x"0e"),
  2822 => (x"86",x"fc",x"0e",x"5d"),
  2823 => (x"6b",x"97",x"4b",x"71"),
  2824 => (x"87",x"e4",x"c0",x"02"),
  2825 => (x"48",x"7e",x"6b",x"97"),
  2826 => (x"a8",x"b7",x"f0",x"c0"),
  2827 => (x"6e",x"87",x"d9",x"04"),
  2828 => (x"b7",x"f9",x"c0",x"48"),
  2829 => (x"87",x"d0",x"01",x"a8"),
  2830 => (x"49",x"6e",x"83",x"c1"),
  2831 => (x"ca",x"89",x"f0",x"c0"),
  2832 => (x"48",x"66",x"d4",x"91"),
  2833 => (x"87",x"c5",x"50",x"71"),
  2834 => (x"eb",x"c4",x"48",x"c0"),
  2835 => (x"02",x"6b",x"97",x"87"),
  2836 => (x"97",x"87",x"e9",x"c0"),
  2837 => (x"c0",x"48",x"7e",x"6b"),
  2838 => (x"04",x"a8",x"b7",x"f0"),
  2839 => (x"48",x"6e",x"87",x"de"),
  2840 => (x"a8",x"b7",x"f9",x"c0"),
  2841 => (x"c1",x"87",x"d5",x"01"),
  2842 => (x"c0",x"49",x"6e",x"83"),
  2843 => (x"66",x"d4",x"89",x"f0"),
  2844 => (x"a1",x"4a",x"bf",x"97"),
  2845 => (x"48",x"66",x"d4",x"49"),
  2846 => (x"87",x"c5",x"50",x"71"),
  2847 => (x"f7",x"c3",x"48",x"c0"),
  2848 => (x"02",x"6b",x"97",x"87"),
  2849 => (x"6b",x"97",x"87",x"cd"),
  2850 => (x"a9",x"fa",x"c0",x"49"),
  2851 => (x"c1",x"87",x"c4",x"05"),
  2852 => (x"c0",x"87",x"c5",x"83"),
  2853 => (x"87",x"e0",x"c3",x"48"),
  2854 => (x"c0",x"02",x"6b",x"97"),
  2855 => (x"6b",x"97",x"87",x"e7"),
  2856 => (x"f0",x"c0",x"48",x"7e"),
  2857 => (x"dc",x"04",x"a8",x"b7"),
  2858 => (x"c0",x"48",x"6e",x"87"),
  2859 => (x"01",x"a8",x"b7",x"f9"),
  2860 => (x"83",x"c1",x"87",x"d3"),
  2861 => (x"f0",x"c0",x"49",x"6e"),
  2862 => (x"d4",x"91",x"ca",x"89"),
  2863 => (x"84",x"c1",x"4c",x"66"),
  2864 => (x"c5",x"7c",x"97",x"71"),
  2865 => (x"c2",x"48",x"c0",x"87"),
  2866 => (x"6b",x"97",x"87",x"ee"),
  2867 => (x"87",x"e4",x"c0",x"02"),
  2868 => (x"48",x"7e",x"6b",x"97"),
  2869 => (x"a8",x"b7",x"f0",x"c0"),
  2870 => (x"6e",x"87",x"d9",x"04"),
  2871 => (x"b7",x"f9",x"c0",x"48"),
  2872 => (x"87",x"d0",x"01",x"a8"),
  2873 => (x"49",x"6e",x"83",x"c1"),
  2874 => (x"97",x"89",x"f0",x"c0"),
  2875 => (x"49",x"a1",x"4a",x"6c"),
  2876 => (x"87",x"c5",x"7c",x"97"),
  2877 => (x"ff",x"c1",x"48",x"c0"),
  2878 => (x"02",x"6b",x"97",x"87"),
  2879 => (x"6b",x"97",x"87",x"cd"),
  2880 => (x"a9",x"fa",x"c0",x"49"),
  2881 => (x"c1",x"87",x"c4",x"05"),
  2882 => (x"c0",x"87",x"c5",x"83"),
  2883 => (x"87",x"e8",x"c1",x"48"),
  2884 => (x"c0",x"02",x"6b",x"97"),
  2885 => (x"6b",x"97",x"87",x"e4"),
  2886 => (x"b7",x"f0",x"c0",x"4a"),
  2887 => (x"87",x"da",x"04",x"aa"),
  2888 => (x"aa",x"b7",x"f9",x"c0"),
  2889 => (x"c1",x"87",x"d3",x"01"),
  2890 => (x"c0",x"49",x"72",x"83"),
  2891 => (x"91",x"ca",x"89",x"f0"),
  2892 => (x"c2",x"4d",x"66",x"d4"),
  2893 => (x"7d",x"97",x"71",x"85"),
  2894 => (x"48",x"c0",x"87",x"c5"),
  2895 => (x"97",x"87",x"f9",x"c0"),
  2896 => (x"e4",x"c0",x"02",x"6b"),
  2897 => (x"7e",x"6b",x"97",x"87"),
  2898 => (x"b7",x"f0",x"c0",x"48"),
  2899 => (x"87",x"d9",x"04",x"a8"),
  2900 => (x"f9",x"c0",x"48",x"6e"),
  2901 => (x"d0",x"01",x"a8",x"b7"),
  2902 => (x"6e",x"83",x"c1",x"87"),
  2903 => (x"89",x"f0",x"c0",x"49"),
  2904 => (x"a1",x"4a",x"6d",x"97"),
  2905 => (x"c4",x"7d",x"97",x"49"),
  2906 => (x"cb",x"48",x"c0",x"87"),
  2907 => (x"02",x"6b",x"97",x"87"),
  2908 => (x"48",x"c0",x"87",x"c4"),
  2909 => (x"48",x"c1",x"87",x"c2"),
  2910 => (x"4d",x"26",x"8e",x"fc"),
  2911 => (x"4b",x"26",x"4c",x"26"),
  2912 => (x"5e",x"0e",x"4f",x"26"),
  2913 => (x"0e",x"5d",x"5c",x"5b"),
  2914 => (x"4d",x"71",x"86",x"f8"),
  2915 => (x"c4",x"4b",x"4c",x"c0"),
  2916 => (x"fd",x"49",x"f8",x"d1"),
  2917 => (x"70",x"87",x"cc",x"fc"),
  2918 => (x"aa",x"b7",x"c0",x"4a"),
  2919 => (x"87",x"f2",x"c2",x"04"),
  2920 => (x"c2",x"02",x"aa",x"ca"),
  2921 => (x"e0",x"c0",x"87",x"ec"),
  2922 => (x"87",x"cf",x"02",x"aa"),
  2923 => (x"ca",x"02",x"aa",x"c9"),
  2924 => (x"02",x"aa",x"cd",x"87"),
  2925 => (x"aa",x"ca",x"87",x"c5"),
  2926 => (x"74",x"87",x"c6",x"05"),
  2927 => (x"d1",x"c2",x"02",x"9c"),
  2928 => (x"aa",x"e2",x"c0",x"87"),
  2929 => (x"74",x"87",x"cc",x"05"),
  2930 => (x"71",x"b9",x"c1",x"49"),
  2931 => (x"9c",x"ff",x"c3",x"4c"),
  2932 => (x"74",x"87",x"fc",x"fe"),
  2933 => (x"e7",x"c1",x"05",x"9c"),
  2934 => (x"b7",x"e1",x"c1",x"87"),
  2935 => (x"87",x"c8",x"04",x"aa"),
  2936 => (x"aa",x"b7",x"fa",x"c1"),
  2937 => (x"87",x"d8",x"c1",x"06"),
  2938 => (x"aa",x"b7",x"c1",x"c1"),
  2939 => (x"c1",x"87",x"c8",x"04"),
  2940 => (x"06",x"aa",x"b7",x"da"),
  2941 => (x"c0",x"87",x"c9",x"c1"),
  2942 => (x"04",x"aa",x"b7",x"f0"),
  2943 => (x"f9",x"c0",x"87",x"c8"),
  2944 => (x"c0",x"06",x"aa",x"b7"),
  2945 => (x"db",x"c1",x"87",x"fa"),
  2946 => (x"f3",x"c0",x"02",x"aa"),
  2947 => (x"aa",x"dd",x"c1",x"87"),
  2948 => (x"87",x"ec",x"c0",x"02"),
  2949 => (x"02",x"aa",x"ed",x"c0"),
  2950 => (x"c1",x"87",x"e5",x"c0"),
  2951 => (x"df",x"02",x"aa",x"df"),
  2952 => (x"aa",x"ec",x"c0",x"87"),
  2953 => (x"c0",x"87",x"d9",x"02"),
  2954 => (x"d3",x"02",x"aa",x"fd"),
  2955 => (x"aa",x"fe",x"c1",x"87"),
  2956 => (x"c0",x"87",x"cd",x"02"),
  2957 => (x"c7",x"02",x"aa",x"fa"),
  2958 => (x"aa",x"ef",x"c0",x"87"),
  2959 => (x"87",x"cf",x"fd",x"05"),
  2960 => (x"ab",x"b7",x"ff",x"c0"),
  2961 => (x"87",x"c7",x"fd",x"03"),
  2962 => (x"c1",x"49",x"a3",x"75"),
  2963 => (x"fc",x"51",x"72",x"83"),
  2964 => (x"a3",x"75",x"87",x"fd"),
  2965 => (x"b7",x"51",x"c0",x"49"),
  2966 => (x"87",x"c4",x"03",x"aa"),
  2967 => (x"87",x"df",x"7e",x"c4"),
  2968 => (x"c7",x"05",x"9b",x"73"),
  2969 => (x"48",x"a6",x"c4",x"87"),
  2970 => (x"87",x"d0",x"78",x"c3"),
  2971 => (x"c4",x"02",x"9c",x"74"),
  2972 => (x"c2",x"7e",x"c1",x"87"),
  2973 => (x"c4",x"7e",x"c0",x"87"),
  2974 => (x"78",x"6e",x"48",x"a6"),
  2975 => (x"6e",x"7e",x"66",x"c4"),
  2976 => (x"26",x"8e",x"f8",x"48"),
  2977 => (x"26",x"4c",x"26",x"4d"),
  2978 => (x"0e",x"4f",x"26",x"4b"),
  2979 => (x"5d",x"5c",x"5b",x"5e"),
  2980 => (x"c4",x"4d",x"71",x"0e"),
  2981 => (x"c0",x"4b",x"c0",x"d1"),
  2982 => (x"49",x"f8",x"c0",x"4a"),
  2983 => (x"87",x"e9",x"c8",x"fd"),
  2984 => (x"d1",x"c4",x"1e",x"75"),
  2985 => (x"eb",x"fd",x"49",x"f8"),
  2986 => (x"86",x"c4",x"87",x"dd"),
  2987 => (x"c5",x"05",x"98",x"70"),
  2988 => (x"c0",x"4c",x"c1",x"87"),
  2989 => (x"49",x"c1",x"87",x"eb"),
  2990 => (x"70",x"87",x"f0",x"c0"),
  2991 => (x"ca",x"05",x"9c",x"4c"),
  2992 => (x"c4",x"d1",x"c4",x"87"),
  2993 => (x"e2",x"c0",x"49",x"bf"),
  2994 => (x"74",x"4c",x"70",x"87"),
  2995 => (x"87",x"cb",x"05",x"9c"),
  2996 => (x"48",x"c0",x"d1",x"c4"),
  2997 => (x"bf",x"d4",x"d1",x"c4"),
  2998 => (x"c4",x"87",x"c6",x"78"),
  2999 => (x"c0",x"48",x"c4",x"d1"),
  3000 => (x"26",x"48",x"74",x"78"),
  3001 => (x"26",x"4c",x"26",x"4d"),
  3002 => (x"0e",x"4f",x"26",x"4b"),
  3003 => (x"5d",x"5c",x"5b",x"5e"),
  3004 => (x"86",x"cc",x"ff",x"0e"),
  3005 => (x"59",x"a6",x"ec",x"c0"),
  3006 => (x"97",x"4c",x"4d",x"c0"),
  3007 => (x"48",x"a6",x"c1",x"7e"),
  3008 => (x"80",x"c0",x"50",x"c0"),
  3009 => (x"c0",x"80",x"c1",x"50"),
  3010 => (x"c0",x"80",x"c4",x"78"),
  3011 => (x"c0",x"80",x"c4",x"78"),
  3012 => (x"c0",x"80",x"c4",x"78"),
  3013 => (x"c0",x"80",x"c4",x"78"),
  3014 => (x"c0",x"d2",x"c4",x"78"),
  3015 => (x"87",x"c5",x"05",x"bf"),
  3016 => (x"d3",x"d0",x"48",x"c1"),
  3017 => (x"f8",x"d1",x"c4",x"87"),
  3018 => (x"d0",x"78",x"c0",x"48"),
  3019 => (x"f4",x"78",x"c0",x"80"),
  3020 => (x"c4",x"d2",x"c4",x"80"),
  3021 => (x"d0",x"c3",x"78",x"bf"),
  3022 => (x"78",x"c0",x"48",x"c0"),
  3023 => (x"48",x"d4",x"d1",x"c4"),
  3024 => (x"cf",x"c3",x"78",x"c0"),
  3025 => (x"f9",x"f8",x"49",x"c0"),
  3026 => (x"58",x"a6",x"dc",x"87"),
  3027 => (x"cd",x"02",x"a8",x"c3"),
  3028 => (x"4b",x"75",x"87",x"d6"),
  3029 => (x"87",x"d8",x"02",x"9b"),
  3030 => (x"c1",x"02",x"8b",x"c1"),
  3031 => (x"02",x"8b",x"87",x"ee"),
  3032 => (x"8b",x"87",x"d3",x"c3"),
  3033 => (x"87",x"f1",x"c6",x"02"),
  3034 => (x"ed",x"c7",x"02",x"8b"),
  3035 => (x"87",x"f8",x"cc",x"87"),
  3036 => (x"cf",x"c3",x"4c",x"c0"),
  3037 => (x"cd",x"c3",x"4a",x"c0"),
  3038 => (x"c3",x"fd",x"49",x"e4"),
  3039 => (x"98",x"70",x"87",x"d1"),
  3040 => (x"c1",x"87",x"c5",x"05"),
  3041 => (x"87",x"e0",x"cc",x"4d"),
  3042 => (x"4a",x"c0",x"cf",x"c3"),
  3043 => (x"49",x"ec",x"cd",x"c3"),
  3044 => (x"87",x"fb",x"c2",x"fd"),
  3045 => (x"c5",x"05",x"98",x"70"),
  3046 => (x"cc",x"4d",x"c2",x"87"),
  3047 => (x"cf",x"c3",x"87",x"ca"),
  3048 => (x"cd",x"c3",x"4a",x"c0"),
  3049 => (x"c2",x"fd",x"49",x"f4"),
  3050 => (x"98",x"70",x"87",x"e5"),
  3051 => (x"87",x"c5",x"c0",x"05"),
  3052 => (x"f3",x"cb",x"4d",x"c3"),
  3053 => (x"c0",x"cf",x"c3",x"87"),
  3054 => (x"fc",x"cd",x"c3",x"4a"),
  3055 => (x"ce",x"c2",x"fd",x"49"),
  3056 => (x"05",x"98",x"70",x"87"),
  3057 => (x"c4",x"87",x"e1",x"cb"),
  3058 => (x"87",x"dc",x"cb",x"4d"),
  3059 => (x"e0",x"c0",x"48",x"74"),
  3060 => (x"98",x"70",x"58",x"a6"),
  3061 => (x"87",x"cb",x"c1",x"05"),
  3062 => (x"c0",x"48",x"a6",x"c8"),
  3063 => (x"66",x"97",x"c2",x"78"),
  3064 => (x"87",x"ca",x"c1",x"05"),
  3065 => (x"bf",x"ec",x"d1",x"c4"),
  3066 => (x"87",x"c7",x"c0",x"02"),
  3067 => (x"50",x"c1",x"80",x"fa"),
  3068 => (x"c3",x"87",x"fb",x"c0"),
  3069 => (x"c4",x"1e",x"c0",x"cf"),
  3070 => (x"fd",x"49",x"e4",x"d1"),
  3071 => (x"c4",x"87",x"c8",x"e6"),
  3072 => (x"02",x"98",x"70",x"86"),
  3073 => (x"c2",x"87",x"c8",x"c0"),
  3074 => (x"50",x"c1",x"48",x"a6"),
  3075 => (x"c4",x"87",x"c3",x"c0"),
  3076 => (x"fe",x"c3",x"7e",x"97"),
  3077 => (x"d1",x"c4",x"1e",x"ec"),
  3078 => (x"ea",x"fd",x"49",x"f8"),
  3079 => (x"86",x"c4",x"87",x"ef"),
  3080 => (x"dc",x"87",x"cb",x"c0"),
  3081 => (x"a8",x"c1",x"48",x"66"),
  3082 => (x"87",x"c2",x"c0",x"05"),
  3083 => (x"84",x"c1",x"4d",x"c0"),
  3084 => (x"c9",x"9c",x"ff",x"c3"),
  3085 => (x"a6",x"d4",x"87",x"f2"),
  3086 => (x"66",x"e0",x"c0",x"48"),
  3087 => (x"c0",x"48",x"74",x"78"),
  3088 => (x"70",x"58",x"a6",x"e0"),
  3089 => (x"fe",x"c0",x"05",x"98"),
  3090 => (x"c0",x"1e",x"ca",x"87"),
  3091 => (x"c0",x"cf",x"c3",x"1e"),
  3092 => (x"ef",x"c4",x"fd",x"49"),
  3093 => (x"70",x"86",x"c8",x"87"),
  3094 => (x"a6",x"e0",x"c0",x"49"),
  3095 => (x"02",x"66",x"dc",x"59"),
  3096 => (x"48",x"87",x"d5",x"c0"),
  3097 => (x"a8",x"b7",x"e3",x"c1"),
  3098 => (x"87",x"cc",x"c0",x"01"),
  3099 => (x"c1",x"49",x"66",x"c4"),
  3100 => (x"a9",x"66",x"dc",x"81"),
  3101 => (x"87",x"c6",x"c0",x"02"),
  3102 => (x"c2",x"7e",x"97",x"c2"),
  3103 => (x"a6",x"c4",x"87",x"d3"),
  3104 => (x"78",x"66",x"dc",x"48"),
  3105 => (x"dc",x"87",x"ca",x"c2"),
  3106 => (x"a8",x"c1",x"48",x"66"),
  3107 => (x"87",x"c1",x"c2",x"05"),
  3108 => (x"4a",x"c0",x"cf",x"c3"),
  3109 => (x"49",x"c4",x"cd",x"c3"),
  3110 => (x"87",x"f3",x"fe",x"fc"),
  3111 => (x"c0",x"05",x"98",x"70"),
  3112 => (x"e0",x"c0",x"87",x"cf"),
  3113 => (x"e4",x"c0",x"48",x"a6"),
  3114 => (x"80",x"c4",x"78",x"f0"),
  3115 => (x"c5",x"c1",x"78",x"c0"),
  3116 => (x"c0",x"cf",x"c3",x"87"),
  3117 => (x"cc",x"cd",x"c3",x"4a"),
  3118 => (x"d2",x"fe",x"fc",x"49"),
  3119 => (x"05",x"98",x"70",x"87"),
  3120 => (x"c0",x"87",x"cf",x"c0"),
  3121 => (x"c0",x"48",x"a6",x"e0"),
  3122 => (x"c4",x"78",x"f0",x"e4"),
  3123 => (x"c0",x"78",x"c1",x"80"),
  3124 => (x"cf",x"c3",x"87",x"e4"),
  3125 => (x"cd",x"c3",x"4a",x"c0"),
  3126 => (x"fd",x"fc",x"49",x"d8"),
  3127 => (x"98",x"70",x"87",x"f1"),
  3128 => (x"87",x"cf",x"c0",x"05"),
  3129 => (x"48",x"a6",x"e0",x"c0"),
  3130 => (x"78",x"c0",x"e0",x"c0"),
  3131 => (x"78",x"c1",x"80",x"c4"),
  3132 => (x"c2",x"87",x"c3",x"c0"),
  3133 => (x"e8",x"c0",x"7e",x"97"),
  3134 => (x"66",x"c4",x"48",x"66"),
  3135 => (x"ce",x"c0",x"05",x"a8"),
  3136 => (x"dc",x"d1",x"c4",x"87"),
  3137 => (x"66",x"e0",x"c0",x"48"),
  3138 => (x"c0",x"80",x"fc",x"78"),
  3139 => (x"c0",x"78",x"66",x"e4"),
  3140 => (x"c3",x"84",x"c1",x"4d"),
  3141 => (x"cf",x"c6",x"9c",x"ff"),
  3142 => (x"a6",x"ec",x"c0",x"87"),
  3143 => (x"c0",x"cf",x"c3",x"1e"),
  3144 => (x"87",x"f0",x"eb",x"49"),
  3145 => (x"98",x"70",x"86",x"c4"),
  3146 => (x"87",x"c6",x"c0",x"05"),
  3147 => (x"c0",x"7e",x"97",x"c2"),
  3148 => (x"ee",x"c0",x"87",x"e3"),
  3149 => (x"1e",x"49",x"66",x"97"),
  3150 => (x"66",x"97",x"f1",x"c0"),
  3151 => (x"f4",x"c0",x"1e",x"49"),
  3152 => (x"ea",x"49",x"66",x"97"),
  3153 => (x"86",x"c8",x"87",x"ec"),
  3154 => (x"d6",x"c2",x"49",x"70"),
  3155 => (x"c8",x"48",x"71",x"81"),
  3156 => (x"a6",x"cc",x"80",x"66"),
  3157 => (x"c5",x"4d",x"c0",x"58"),
  3158 => (x"48",x"74",x"87",x"ce"),
  3159 => (x"58",x"a6",x"e0",x"c0"),
  3160 => (x"c0",x"05",x"98",x"70"),
  3161 => (x"1e",x"ca",x"87",x"d7"),
  3162 => (x"cf",x"c3",x"1e",x"c0"),
  3163 => (x"c0",x"fd",x"49",x"c0"),
  3164 => (x"86",x"c8",x"87",x"d2"),
  3165 => (x"a6",x"c5",x"49",x"70"),
  3166 => (x"e6",x"c4",x"59",x"97"),
  3167 => (x"48",x"66",x"dc",x"87"),
  3168 => (x"c4",x"05",x"a8",x"c1"),
  3169 => (x"ec",x"c0",x"87",x"dd"),
  3170 => (x"cf",x"c3",x"1e",x"a6"),
  3171 => (x"c3",x"ea",x"49",x"c0"),
  3172 => (x"70",x"86",x"c4",x"87"),
  3173 => (x"c6",x"c0",x"05",x"98"),
  3174 => (x"7e",x"97",x"c2",x"87"),
  3175 => (x"c0",x"87",x"c2",x"c4"),
  3176 => (x"49",x"66",x"97",x"ee"),
  3177 => (x"97",x"f1",x"c0",x"1e"),
  3178 => (x"c0",x"1e",x"49",x"66"),
  3179 => (x"49",x"66",x"97",x"f4"),
  3180 => (x"c8",x"87",x"ff",x"e8"),
  3181 => (x"a6",x"e0",x"c0",x"86"),
  3182 => (x"66",x"97",x"c1",x"58"),
  3183 => (x"a6",x"f4",x"c0",x"48"),
  3184 => (x"05",x"98",x"70",x"58"),
  3185 => (x"c0",x"87",x"e7",x"c0"),
  3186 => (x"c1",x"49",x"66",x"e8"),
  3187 => (x"a9",x"66",x"c4",x"81"),
  3188 => (x"87",x"cd",x"c3",x"05"),
  3189 => (x"bf",x"d4",x"d1",x"c4"),
  3190 => (x"87",x"c5",x"c3",x"05"),
  3191 => (x"c2",x"49",x"66",x"dc"),
  3192 => (x"48",x"71",x"81",x"d6"),
  3193 => (x"c4",x"80",x"66",x"c8"),
  3194 => (x"c2",x"58",x"d8",x"d1"),
  3195 => (x"f0",x"c0",x"87",x"f3"),
  3196 => (x"a8",x"c1",x"48",x"66"),
  3197 => (x"87",x"e9",x"c2",x"05"),
  3198 => (x"c0",x"48",x"66",x"c4"),
  3199 => (x"05",x"a8",x"66",x"e8"),
  3200 => (x"dc",x"87",x"cf",x"c0"),
  3201 => (x"d6",x"c2",x"49",x"66"),
  3202 => (x"c8",x"48",x"71",x"81"),
  3203 => (x"d1",x"c4",x"80",x"66"),
  3204 => (x"66",x"c4",x"58",x"d4"),
  3205 => (x"a8",x"b7",x"c1",x"48"),
  3206 => (x"87",x"dd",x"c1",x"06"),
  3207 => (x"cc",x"48",x"66",x"dc"),
  3208 => (x"f4",x"c0",x"88",x"66"),
  3209 => (x"66",x"c4",x"58",x"a6"),
  3210 => (x"66",x"e8",x"c0",x"48"),
  3211 => (x"d0",x"c0",x"05",x"a8"),
  3212 => (x"66",x"f0",x"c0",x"87"),
  3213 => (x"91",x"66",x"d4",x"49"),
  3214 => (x"66",x"d0",x"48",x"71"),
  3215 => (x"d0",x"d1",x"c4",x"80"),
  3216 => (x"66",x"e8",x"c0",x"58"),
  3217 => (x"c4",x"81",x"c1",x"49"),
  3218 => (x"c0",x"05",x"a9",x"66"),
  3219 => (x"d1",x"c4",x"87",x"d9"),
  3220 => (x"c0",x"05",x"bf",x"d4"),
  3221 => (x"66",x"dc",x"87",x"d1"),
  3222 => (x"81",x"d6",x"c2",x"49"),
  3223 => (x"71",x"81",x"66",x"c8"),
  3224 => (x"c4",x"88",x"c1",x"48"),
  3225 => (x"c0",x"58",x"d8",x"d1"),
  3226 => (x"d4",x"49",x"66",x"f0"),
  3227 => (x"48",x"71",x"91",x"66"),
  3228 => (x"d4",x"80",x"66",x"d0"),
  3229 => (x"e2",x"c0",x"58",x"a6"),
  3230 => (x"49",x"66",x"dc",x"87"),
  3231 => (x"d4",x"81",x"d6",x"c2"),
  3232 => (x"48",x"71",x"91",x"66"),
  3233 => (x"d4",x"80",x"66",x"d0"),
  3234 => (x"e8",x"c0",x"58",x"a6"),
  3235 => (x"a8",x"c1",x"48",x"66"),
  3236 => (x"87",x"c7",x"c0",x"05"),
  3237 => (x"48",x"cc",x"d1",x"c4"),
  3238 => (x"cc",x"78",x"66",x"d0"),
  3239 => (x"66",x"dc",x"48",x"a6"),
  3240 => (x"c1",x"4d",x"c0",x"78"),
  3241 => (x"9c",x"ff",x"c3",x"84"),
  3242 => (x"c4",x"48",x"66",x"d8"),
  3243 => (x"c6",x"c0",x"02",x"a8"),
  3244 => (x"02",x"6e",x"97",x"87"),
  3245 => (x"c2",x"87",x"cb",x"f2"),
  3246 => (x"c0",x"05",x"66",x"97"),
  3247 => (x"97",x"c4",x"87",x"c6"),
  3248 => (x"87",x"f6",x"c0",x"7e"),
  3249 => (x"c0",x"48",x"66",x"c4"),
  3250 => (x"05",x"a8",x"66",x"e8"),
  3251 => (x"c4",x"87",x"eb",x"c0"),
  3252 => (x"4a",x"bf",x"cc",x"d1"),
  3253 => (x"bf",x"ec",x"d1",x"c4"),
  3254 => (x"70",x"88",x"72",x"48"),
  3255 => (x"dc",x"d1",x"c4",x"4a"),
  3256 => (x"1e",x"72",x"49",x"bf"),
  3257 => (x"fc",x"4a",x"09",x"72"),
  3258 => (x"70",x"87",x"e7",x"fc"),
  3259 => (x"c4",x"4a",x"26",x"49"),
  3260 => (x"48",x"bf",x"d0",x"d1"),
  3261 => (x"d1",x"c4",x"80",x"71"),
  3262 => (x"66",x"c4",x"58",x"d8"),
  3263 => (x"66",x"e8",x"c0",x"48"),
  3264 => (x"c0",x"03",x"a8",x"b7"),
  3265 => (x"97",x"c4",x"87",x"c3"),
  3266 => (x"02",x"6e",x"97",x"7e"),
  3267 => (x"c4",x"87",x"c9",x"c0"),
  3268 => (x"c0",x"48",x"c4",x"d1"),
  3269 => (x"87",x"c7",x"c0",x"78"),
  3270 => (x"48",x"c4",x"d1",x"c4"),
  3271 => (x"c0",x"78",x"66",x"c4"),
  3272 => (x"c4",x"1e",x"a6",x"ec"),
  3273 => (x"49",x"bf",x"d0",x"d1"),
  3274 => (x"c4",x"87",x"fd",x"e1"),
  3275 => (x"e0",x"d1",x"c4",x"86"),
  3276 => (x"66",x"e8",x"c0",x"48"),
  3277 => (x"48",x"6e",x"97",x"78"),
  3278 => (x"26",x"8e",x"cc",x"ff"),
  3279 => (x"26",x"4c",x"26",x"4d"),
  3280 => (x"00",x"4f",x"26",x"4b"),
  3281 => (x"49",x"44",x"55",x"41"),
  3282 => (x"00",x"00",x"00",x"4f"),
  3283 => (x"45",x"44",x"4f",x"4d"),
  3284 => (x"33",x"32",x"2f",x"31"),
  3285 => (x"00",x"00",x"32",x"35"),
  3286 => (x"45",x"44",x"4f",x"4d"),
  3287 => (x"30",x"32",x"2f",x"31"),
  3288 => (x"00",x"00",x"38",x"34"),
  3289 => (x"45",x"4c",x"49",x"46"),
  3290 => (x"00",x"00",x"00",x"00"),
  3291 => (x"43",x"41",x"52",x"54"),
  3292 => (x"00",x"00",x"00",x"4b"),
  3293 => (x"47",x"45",x"52",x"50"),
  3294 => (x"00",x"00",x"50",x"41"),
  3295 => (x"45",x"44",x"4e",x"49"),
  3296 => (x"5e",x"0e",x"00",x"58"),
  3297 => (x"71",x"0e",x"5c",x"5b"),
  3298 => (x"c4",x"4b",x"c1",x"4c"),
  3299 => (x"b7",x"bf",x"d0",x"d1"),
  3300 => (x"87",x"d0",x"04",x"ac"),
  3301 => (x"bf",x"d4",x"d1",x"c4"),
  3302 => (x"c7",x"01",x"ac",x"b7"),
  3303 => (x"e0",x"d1",x"c4",x"87"),
  3304 => (x"87",x"d3",x"48",x"bf"),
  3305 => (x"c2",x"ed",x"49",x"73"),
  3306 => (x"c4",x"83",x"c1",x"87"),
  3307 => (x"b7",x"bf",x"c4",x"d1"),
  3308 => (x"d6",x"ff",x"06",x"ab"),
  3309 => (x"26",x"48",x"ff",x"87"),
  3310 => (x"26",x"4b",x"26",x"4c"),
  3311 => (x"00",x"00",x"00",x"4f"),
  3312 => (x"00",x"00",x"00",x"00"),
  3313 => (x"00",x"00",x"00",x"00"),
  3314 => (x"00",x"00",x"00",x"00"),
  3315 => (x"00",x"00",x"00",x"00"),
  3316 => (x"00",x"00",x"00",x"00"),
  3317 => (x"00",x"00",x"00",x"00"),
  3318 => (x"00",x"00",x"00",x"00"),
  3319 => (x"00",x"00",x"00",x"00"),
  3320 => (x"00",x"00",x"00",x"00"),
  3321 => (x"00",x"00",x"00",x"00"),
  3322 => (x"00",x"00",x"00",x"00"),
  3323 => (x"00",x"00",x"00",x"00"),
  3324 => (x"00",x"00",x"00",x"00"),
  3325 => (x"00",x"00",x"00",x"00"),
  3326 => (x"00",x"00",x"00",x"00"),
  3327 => (x"00",x"00",x"00",x"00"),
  3328 => (x"00",x"00",x"00",x"00"),
  3329 => (x"71",x"1e",x"73",x"1e"),
  3330 => (x"72",x"1e",x"4a",x"4b"),
  3331 => (x"fc",x"4a",x"ca",x"49"),
  3332 => (x"70",x"87",x"f3",x"f8"),
  3333 => (x"d0",x"4a",x"26",x"49"),
  3334 => (x"72",x"1e",x"71",x"91"),
  3335 => (x"fc",x"4a",x"ca",x"49"),
  3336 => (x"71",x"87",x"e3",x"f8"),
  3337 => (x"72",x"49",x"26",x"4a"),
  3338 => (x"ff",x"c3",x"49",x"a1"),
  3339 => (x"26",x"48",x"71",x"99"),
  3340 => (x"1e",x"4f",x"26",x"4b"),
  3341 => (x"4b",x"71",x"1e",x"73"),
  3342 => (x"b7",x"c4",x"49",x"4a"),
  3343 => (x"cf",x"91",x"ca",x"29"),
  3344 => (x"49",x"a1",x"72",x"9a"),
  3345 => (x"71",x"99",x"ff",x"c3"),
  3346 => (x"26",x"4b",x"26",x"48"),
  3347 => (x"1e",x"73",x"1e",x"4f"),
  3348 => (x"ff",x"49",x"4a",x"71"),
  3349 => (x"49",x"70",x"87",x"dd"),
  3350 => (x"c2",x"05",x"9b",x"4b"),
  3351 => (x"c4",x"4b",x"c1",x"87"),
  3352 => (x"b7",x"bf",x"c4",x"d1"),
  3353 => (x"87",x"c1",x"06",x"ab"),
  3354 => (x"e9",x"49",x"73",x"4b"),
  3355 => (x"48",x"73",x"87",x"fd"),
  3356 => (x"4f",x"26",x"4b",x"26"),
  3357 => (x"c0",x"f7",x"c4",x"1e"),
  3358 => (x"f6",x"c4",x"59",x"97"),
  3359 => (x"66",x"c4",x"48",x"fd"),
  3360 => (x"50",x"66",x"c8",x"50"),
  3361 => (x"26",x"50",x"66",x"cc"),
  3362 => (x"1e",x"73",x"1e",x"4f"),
  3363 => (x"d0",x"ff",x"4b",x"71"),
  3364 => (x"78",x"c5",x"c8",x"48"),
  3365 => (x"c1",x"48",x"d4",x"ff"),
  3366 => (x"49",x"73",x"78",x"e1"),
  3367 => (x"2a",x"b7",x"c8",x"4a"),
  3368 => (x"ff",x"c3",x"78",x"72"),
  3369 => (x"ff",x"78",x"71",x"99"),
  3370 => (x"78",x"c4",x"48",x"d0"),
  3371 => (x"4f",x"26",x"4b",x"26"),
  3372 => (x"fe",x"f7",x"c4",x"1e"),
  3373 => (x"f7",x"c4",x"59",x"9f"),
  3374 => (x"78",x"c1",x"48",x"cc"),
  3375 => (x"5e",x"0e",x"4f",x"26"),
  3376 => (x"71",x"0e",x"5c",x"5b"),
  3377 => (x"48",x"d0",x"ff",x"4c"),
  3378 => (x"ff",x"78",x"c5",x"c8"),
  3379 => (x"e4",x"c1",x"48",x"d4"),
  3380 => (x"49",x"66",x"cc",x"78"),
  3381 => (x"9a",x"ff",x"c3",x"4a"),
  3382 => (x"66",x"cc",x"78",x"72"),
  3383 => (x"c3",x"2a",x"c8",x"4a"),
  3384 => (x"66",x"d0",x"9a",x"ff"),
  3385 => (x"73",x"33",x"c7",x"4b"),
  3386 => (x"71",x"78",x"72",x"b2"),
  3387 => (x"fc",x"49",x"74",x"1e"),
  3388 => (x"ff",x"87",x"c4",x"f6"),
  3389 => (x"78",x"c4",x"48",x"d0"),
  3390 => (x"4c",x"26",x"8e",x"fc"),
  3391 => (x"4f",x"26",x"4b",x"26"),
  3392 => (x"c0",x"1e",x"73",x"1e"),
  3393 => (x"c4",x"4b",x"c0",x"e0"),
  3394 => (x"02",x"bf",x"d8",x"d1"),
  3395 => (x"c4",x"87",x"e7",x"c1"),
  3396 => (x"48",x"bf",x"d8",x"f7"),
  3397 => (x"04",x"a8",x"b7",x"c0"),
  3398 => (x"c4",x"87",x"db",x"c1"),
  3399 => (x"ab",x"bf",x"dc",x"d1"),
  3400 => (x"c4",x"87",x"d3",x"02"),
  3401 => (x"49",x"bf",x"f4",x"d1"),
  3402 => (x"1e",x"71",x"81",x"d0"),
  3403 => (x"49",x"e4",x"d1",x"c4"),
  3404 => (x"87",x"e9",x"d7",x"fd"),
  3405 => (x"1e",x"73",x"86",x"c4"),
  3406 => (x"1e",x"cc",x"d2",x"c4"),
  3407 => (x"49",x"e4",x"d1",x"c4"),
  3408 => (x"87",x"c2",x"d9",x"fd"),
  3409 => (x"d1",x"c4",x"86",x"c8"),
  3410 => (x"02",x"ab",x"bf",x"dc"),
  3411 => (x"c0",x"49",x"87",x"d6"),
  3412 => (x"c4",x"89",x"d0",x"e0"),
  3413 => (x"81",x"bf",x"f4",x"d1"),
  3414 => (x"d1",x"c4",x"1e",x"71"),
  3415 => (x"d6",x"fd",x"49",x"e4"),
  3416 => (x"86",x"c4",x"87",x"fb"),
  3417 => (x"1e",x"49",x"66",x"c8"),
  3418 => (x"d2",x"c4",x"1e",x"73"),
  3419 => (x"cd",x"fd",x"49",x"cc"),
  3420 => (x"c0",x"86",x"c8",x"87"),
  3421 => (x"e4",x"c0",x"87",x"e1"),
  3422 => (x"d2",x"c4",x"1e",x"f0"),
  3423 => (x"d1",x"c4",x"1e",x"cc"),
  3424 => (x"d8",x"fd",x"49",x"e4"),
  3425 => (x"66",x"d0",x"87",x"c0"),
  3426 => (x"e4",x"c0",x"1e",x"49"),
  3427 => (x"d2",x"c4",x"1e",x"f0"),
  3428 => (x"e9",x"fc",x"49",x"cc"),
  3429 => (x"26",x"86",x"d0",x"87"),
  3430 => (x"1e",x"4f",x"26",x"4b"),
  3431 => (x"bf",x"ec",x"d1",x"c4"),
  3432 => (x"c4",x"87",x"db",x"05"),
  3433 => (x"c1",x"48",x"c4",x"f7"),
  3434 => (x"1e",x"1e",x"c0",x"50"),
  3435 => (x"49",x"c2",x"1e",x"cb"),
  3436 => (x"cc",x"87",x"c1",x"fb"),
  3437 => (x"fb",x"49",x"c1",x"86"),
  3438 => (x"48",x"c0",x"87",x"cf"),
  3439 => (x"48",x"c1",x"87",x"c2"),
  3440 => (x"5e",x"0e",x"4f",x"26"),
  3441 => (x"c0",x"0e",x"5c",x"5b"),
  3442 => (x"c4",x"4c",x"f0",x"e4"),
  3443 => (x"48",x"bf",x"c0",x"f7"),
  3444 => (x"c0",x"06",x"a8",x"c0"),
  3445 => (x"fb",x"c3",x"87",x"e9"),
  3446 => (x"c0",x"49",x"bf",x"cc"),
  3447 => (x"70",x"87",x"fd",x"e3"),
  3448 => (x"df",x"c7",x"02",x"98"),
  3449 => (x"c0",x"49",x"cd",x"87"),
  3450 => (x"70",x"87",x"e5",x"e3"),
  3451 => (x"d0",x"fb",x"c3",x"49"),
  3452 => (x"c0",x"f7",x"c4",x"59"),
  3453 => (x"88",x"c1",x"48",x"bf"),
  3454 => (x"58",x"c4",x"f7",x"c4"),
  3455 => (x"c4",x"87",x"c5",x"c7"),
  3456 => (x"bf",x"97",x"c4",x"f7"),
  3457 => (x"05",x"aa",x"c2",x"4a"),
  3458 => (x"c4",x"87",x"ca",x"c3"),
  3459 => (x"48",x"bf",x"d4",x"f7"),
  3460 => (x"bf",x"c4",x"d1",x"c4"),
  3461 => (x"c9",x"06",x"a8",x"b7"),
  3462 => (x"c4",x"f7",x"c4",x"87"),
  3463 => (x"c6",x"50",x"c0",x"48"),
  3464 => (x"f7",x"c4",x"87",x"e2"),
  3465 => (x"02",x"bf",x"97",x"d1"),
  3466 => (x"c4",x"87",x"d9",x"c6"),
  3467 => (x"05",x"bf",x"ec",x"d1"),
  3468 => (x"f7",x"c4",x"87",x"da"),
  3469 => (x"50",x"c1",x"48",x"c4"),
  3470 => (x"cb",x"1e",x"1e",x"c0"),
  3471 => (x"f8",x"49",x"c2",x"1e"),
  3472 => (x"86",x"cc",x"87",x"f2"),
  3473 => (x"e7",x"f9",x"49",x"c1"),
  3474 => (x"87",x"f8",x"c5",x"87"),
  3475 => (x"48",x"d1",x"f7",x"c4"),
  3476 => (x"d1",x"c4",x"50",x"c0"),
  3477 => (x"cd",x"02",x"bf",x"d8"),
  3478 => (x"c0",x"1e",x"c1",x"87"),
  3479 => (x"fa",x"49",x"c0",x"e0"),
  3480 => (x"86",x"c4",x"87",x"de"),
  3481 => (x"f7",x"c4",x"87",x"d5"),
  3482 => (x"c4",x"48",x"bf",x"d8"),
  3483 => (x"b7",x"bf",x"d0",x"d1"),
  3484 => (x"c6",x"c0",x"04",x"a8"),
  3485 => (x"c5",x"f7",x"c4",x"87"),
  3486 => (x"c4",x"50",x"c0",x"48"),
  3487 => (x"48",x"bf",x"dc",x"f7"),
  3488 => (x"f7",x"c4",x"88",x"c1"),
  3489 => (x"98",x"70",x"58",x"e0"),
  3490 => (x"87",x"cb",x"c0",x"05"),
  3491 => (x"df",x"f8",x"49",x"c0"),
  3492 => (x"c4",x"f7",x"c4",x"87"),
  3493 => (x"c4",x"50",x"c0",x"48"),
  3494 => (x"48",x"bf",x"d8",x"f7"),
  3495 => (x"f7",x"c4",x"80",x"c1"),
  3496 => (x"d1",x"c4",x"58",x"dc"),
  3497 => (x"a8",x"b7",x"bf",x"d4"),
  3498 => (x"87",x"d8",x"c4",x"04"),
  3499 => (x"bf",x"d4",x"f7",x"c4"),
  3500 => (x"c4",x"80",x"c1",x"48"),
  3501 => (x"70",x"58",x"d8",x"f7"),
  3502 => (x"87",x"ef",x"e0",x"49"),
  3503 => (x"48",x"c5",x"f7",x"c4"),
  3504 => (x"d1",x"c4",x"50",x"c1"),
  3505 => (x"1e",x"49",x"bf",x"cc"),
  3506 => (x"49",x"e4",x"d1",x"c4"),
  3507 => (x"87",x"cd",x"d1",x"fd"),
  3508 => (x"ef",x"c3",x"86",x"c4"),
  3509 => (x"05",x"aa",x"c3",x"87"),
  3510 => (x"c4",x"87",x"e9",x"c3"),
  3511 => (x"05",x"bf",x"ec",x"d1"),
  3512 => (x"c4",x"87",x"da",x"c0"),
  3513 => (x"c1",x"48",x"c4",x"f7"),
  3514 => (x"1e",x"1e",x"c0",x"50"),
  3515 => (x"49",x"c2",x"1e",x"cb"),
  3516 => (x"cc",x"87",x"c1",x"f6"),
  3517 => (x"f6",x"49",x"c1",x"86"),
  3518 => (x"c7",x"c3",x"87",x"f6"),
  3519 => (x"d8",x"f7",x"c4",x"87"),
  3520 => (x"fd",x"f1",x"49",x"bf"),
  3521 => (x"d8",x"f7",x"c4",x"87"),
  3522 => (x"d2",x"f7",x"c4",x"58"),
  3523 => (x"c1",x"05",x"bf",x"97"),
  3524 => (x"4b",x"c0",x"87",x"d1"),
  3525 => (x"bf",x"f4",x"f7",x"c4"),
  3526 => (x"a8",x"b7",x"c0",x"48"),
  3527 => (x"87",x"c3",x"c1",x"04"),
  3528 => (x"bf",x"d8",x"d1",x"c4"),
  3529 => (x"87",x"e4",x"c0",x"05"),
  3530 => (x"bf",x"d8",x"f7",x"c4"),
  3531 => (x"d0",x"d1",x"c4",x"49"),
  3532 => (x"91",x"74",x"89",x"bf"),
  3533 => (x"bf",x"cc",x"d1",x"c4"),
  3534 => (x"c4",x"1e",x"71",x"81"),
  3535 => (x"fd",x"49",x"e4",x"d1"),
  3536 => (x"c0",x"87",x"da",x"cf"),
  3537 => (x"f6",x"49",x"74",x"1e"),
  3538 => (x"86",x"c8",x"87",x"f6"),
  3539 => (x"bf",x"d8",x"f7",x"c4"),
  3540 => (x"c4",x"80",x"c1",x"48"),
  3541 => (x"c1",x"58",x"dc",x"f7"),
  3542 => (x"f4",x"f7",x"c4",x"83"),
  3543 => (x"06",x"ab",x"b7",x"bf"),
  3544 => (x"c4",x"87",x"fd",x"fe"),
  3545 => (x"c0",x"48",x"f4",x"f7"),
  3546 => (x"d8",x"f7",x"c4",x"78"),
  3547 => (x"f7",x"c4",x"48",x"bf"),
  3548 => (x"a8",x"b7",x"bf",x"f0"),
  3549 => (x"87",x"d7",x"c0",x"03"),
  3550 => (x"bf",x"d8",x"d1",x"c4"),
  3551 => (x"87",x"cf",x"c0",x"05"),
  3552 => (x"bf",x"d4",x"f7",x"c4"),
  3553 => (x"c4",x"d1",x"c4",x"48"),
  3554 => (x"06",x"a8",x"b7",x"bf"),
  3555 => (x"c4",x"87",x"f5",x"c0"),
  3556 => (x"bf",x"97",x"f8",x"f7"),
  3557 => (x"05",x"a9",x"c1",x"49"),
  3558 => (x"c4",x"87",x"d2",x"c0"),
  3559 => (x"c4",x"48",x"d8",x"f7"),
  3560 => (x"78",x"bf",x"ec",x"f7"),
  3561 => (x"48",x"c0",x"f7",x"c4"),
  3562 => (x"c6",x"c0",x"78",x"c2"),
  3563 => (x"c4",x"f7",x"c4",x"87"),
  3564 => (x"c4",x"50",x"c0",x"48"),
  3565 => (x"bf",x"97",x"f8",x"f7"),
  3566 => (x"05",x"a9",x"c2",x"49"),
  3567 => (x"c0",x"87",x"c5",x"c0"),
  3568 => (x"87",x"ec",x"f3",x"49"),
  3569 => (x"4b",x"26",x"4c",x"26"),
  3570 => (x"5e",x"0e",x"4f",x"26"),
  3571 => (x"0e",x"5d",x"5c",x"5b"),
  3572 => (x"76",x"86",x"c4",x"ff"),
  3573 => (x"c0",x"4a",x"c0",x"4b"),
  3574 => (x"e3",x"fc",x"49",x"e0"),
  3575 => (x"d0",x"ff",x"87",x"eb"),
  3576 => (x"78",x"c5",x"c8",x"48"),
  3577 => (x"c1",x"48",x"d4",x"ff"),
  3578 => (x"4d",x"c0",x"78",x"e2"),
  3579 => (x"7c",x"c0",x"4c",x"70"),
  3580 => (x"49",x"a6",x"e0",x"c0"),
  3581 => (x"51",x"6c",x"81",x"75"),
  3582 => (x"b7",x"cc",x"85",x"c1"),
  3583 => (x"87",x"ee",x"04",x"ad"),
  3584 => (x"c4",x"48",x"d0",x"ff"),
  3585 => (x"97",x"e0",x"c0",x"78"),
  3586 => (x"02",x"9c",x"4c",x"66"),
  3587 => (x"c3",x"87",x"f3",x"c0"),
  3588 => (x"fe",x"c0",x"02",x"8c"),
  3589 => (x"02",x"8c",x"c5",x"87"),
  3590 => (x"cd",x"87",x"e7",x"c6"),
  3591 => (x"f3",x"c8",x"02",x"8c"),
  3592 => (x"8c",x"c3",x"c3",x"87"),
  3593 => (x"87",x"c5",x"c9",x"02"),
  3594 => (x"cc",x"02",x"8c",x"c1"),
  3595 => (x"02",x"8c",x"87",x"e9"),
  3596 => (x"c3",x"87",x"ee",x"d0"),
  3597 => (x"ff",x"d0",x"02",x"8c"),
  3598 => (x"02",x"8c",x"c1",x"87"),
  3599 => (x"d4",x"87",x"f8",x"c1"),
  3600 => (x"d6",x"f5",x"87",x"f1"),
  3601 => (x"02",x"98",x"70",x"87"),
  3602 => (x"c0",x"87",x"c2",x"d5"),
  3603 => (x"87",x"f9",x"f0",x"49"),
  3604 => (x"d2",x"87",x"fa",x"d4"),
  3605 => (x"a6",x"c1",x"7e",x"97"),
  3606 => (x"50",x"c0",x"c2",x"48"),
  3607 => (x"c1",x"50",x"f0",x"c1"),
  3608 => (x"fc",x"f6",x"c4",x"80"),
  3609 => (x"c4",x"50",x"bf",x"97"),
  3610 => (x"c4",x"50",x"ca",x"80"),
  3611 => (x"fd",x"f6",x"c4",x"80"),
  3612 => (x"c4",x"50",x"bf",x"97"),
  3613 => (x"bf",x"97",x"fe",x"f6"),
  3614 => (x"ff",x"f6",x"c4",x"50"),
  3615 => (x"c4",x"50",x"bf",x"97"),
  3616 => (x"c0",x"48",x"ff",x"f6"),
  3617 => (x"fe",x"f6",x"c4",x"50"),
  3618 => (x"ff",x"f6",x"c4",x"48"),
  3619 => (x"c4",x"50",x"bf",x"97"),
  3620 => (x"c4",x"48",x"fd",x"f6"),
  3621 => (x"bf",x"97",x"fe",x"f6"),
  3622 => (x"fc",x"f6",x"c4",x"50"),
  3623 => (x"fd",x"f6",x"c4",x"48"),
  3624 => (x"c1",x"50",x"bf",x"97"),
  3625 => (x"ca",x"1e",x"d2",x"1e"),
  3626 => (x"d1",x"f0",x"49",x"a6"),
  3627 => (x"c0",x"86",x"c8",x"87"),
  3628 => (x"87",x"d5",x"ef",x"49"),
  3629 => (x"f3",x"87",x"d6",x"d3"),
  3630 => (x"98",x"70",x"87",x"e1"),
  3631 => (x"87",x"cd",x"d3",x"02"),
  3632 => (x"66",x"97",x"e1",x"c0"),
  3633 => (x"a6",x"f0",x"c0",x"48"),
  3634 => (x"02",x"98",x"70",x"58"),
  3635 => (x"c1",x"48",x"87",x"da"),
  3636 => (x"a6",x"f0",x"c0",x"88"),
  3637 => (x"02",x"98",x"70",x"58"),
  3638 => (x"48",x"87",x"ed",x"c0"),
  3639 => (x"f0",x"c0",x"88",x"c1"),
  3640 => (x"98",x"70",x"58",x"a6"),
  3641 => (x"87",x"ec",x"c1",x"02"),
  3642 => (x"c1",x"7e",x"97",x"c2"),
  3643 => (x"c0",x"c2",x"48",x"a6"),
  3644 => (x"c4",x"50",x"c1",x"50"),
  3645 => (x"49",x"bf",x"c4",x"d1"),
  3646 => (x"c3",x"87",x"c9",x"ec"),
  3647 => (x"c0",x"50",x"08",x"a6"),
  3648 => (x"c2",x"48",x"a6",x"ec"),
  3649 => (x"87",x"e4",x"c2",x"78"),
  3650 => (x"bf",x"c0",x"d1",x"c4"),
  3651 => (x"81",x"d6",x"c2",x"49"),
  3652 => (x"1e",x"a6",x"f0",x"c0"),
  3653 => (x"cf",x"ca",x"ff",x"71"),
  3654 => (x"97",x"86",x"c4",x"87"),
  3655 => (x"48",x"a6",x"c1",x"7e"),
  3656 => (x"c0",x"50",x"c0",x"c2"),
  3657 => (x"49",x"66",x"97",x"f0"),
  3658 => (x"c2",x"87",x"d9",x"eb"),
  3659 => (x"c0",x"50",x"08",x"a6"),
  3660 => (x"49",x"66",x"97",x"f1"),
  3661 => (x"c3",x"87",x"cd",x"eb"),
  3662 => (x"c0",x"50",x"08",x"a6"),
  3663 => (x"49",x"66",x"97",x"f2"),
  3664 => (x"c4",x"87",x"c1",x"eb"),
  3665 => (x"c5",x"50",x"08",x"a6"),
  3666 => (x"50",x"c0",x"48",x"a6"),
  3667 => (x"c4",x"80",x"e6",x"c0"),
  3668 => (x"87",x"d8",x"c1",x"78"),
  3669 => (x"66",x"97",x"e2",x"c0"),
  3670 => (x"87",x"f1",x"eb",x"49"),
  3671 => (x"bf",x"d0",x"d1",x"c4"),
  3672 => (x"81",x"d6",x"c2",x"49"),
  3673 => (x"1e",x"a6",x"f0",x"c0"),
  3674 => (x"fb",x"c8",x"ff",x"71"),
  3675 => (x"97",x"86",x"c4",x"87"),
  3676 => (x"48",x"a6",x"c1",x"7e"),
  3677 => (x"c0",x"50",x"c0",x"c2"),
  3678 => (x"49",x"66",x"97",x"f0"),
  3679 => (x"c2",x"87",x"c5",x"ea"),
  3680 => (x"c0",x"50",x"08",x"a6"),
  3681 => (x"49",x"66",x"97",x"f1"),
  3682 => (x"c3",x"87",x"f9",x"e9"),
  3683 => (x"c0",x"50",x"08",x"a6"),
  3684 => (x"49",x"66",x"97",x"f2"),
  3685 => (x"c4",x"87",x"ed",x"e9"),
  3686 => (x"c4",x"50",x"08",x"a6"),
  3687 => (x"49",x"bf",x"d8",x"d1"),
  3688 => (x"a6",x"c9",x"31",x"c2"),
  3689 => (x"c0",x"48",x"59",x"97"),
  3690 => (x"78",x"c4",x"80",x"e7"),
  3691 => (x"f0",x"c0",x"1e",x"c1"),
  3692 => (x"a6",x"ca",x"1e",x"66"),
  3693 => (x"87",x"c6",x"ec",x"49"),
  3694 => (x"49",x"c0",x"86",x"c8"),
  3695 => (x"cf",x"87",x"ca",x"eb"),
  3696 => (x"d6",x"ef",x"87",x"cb"),
  3697 => (x"02",x"98",x"70",x"87"),
  3698 => (x"c0",x"87",x"c2",x"cf"),
  3699 => (x"49",x"66",x"97",x"e1"),
  3700 => (x"e2",x"c0",x"31",x"d0"),
  3701 => (x"c8",x"4a",x"66",x"97"),
  3702 => (x"c0",x"b1",x"72",x"32"),
  3703 => (x"4a",x"66",x"97",x"e3"),
  3704 => (x"c7",x"48",x"71",x"b1"),
  3705 => (x"98",x"ff",x"ff",x"ff"),
  3706 => (x"58",x"a6",x"f0",x"c0"),
  3707 => (x"66",x"97",x"e4",x"c0"),
  3708 => (x"87",x"c8",x"c0",x"02"),
  3709 => (x"a6",x"f8",x"c0",x"48"),
  3710 => (x"87",x"c7",x"c0",x"58"),
  3711 => (x"48",x"a6",x"f4",x"c0"),
  3712 => (x"c0",x"78",x"c0",x"c4"),
  3713 => (x"e5",x"49",x"66",x"ec"),
  3714 => (x"f7",x"c4",x"87",x"f8"),
  3715 => (x"f7",x"c4",x"58",x"d8"),
  3716 => (x"78",x"c0",x"48",x"c0"),
  3717 => (x"48",x"d8",x"f7",x"c4"),
  3718 => (x"40",x"66",x"ec",x"c0"),
  3719 => (x"78",x"66",x"f4",x"c0"),
  3720 => (x"49",x"66",x"ec",x"c0"),
  3721 => (x"bf",x"d0",x"d1",x"c4"),
  3722 => (x"dc",x"d1",x"c4",x"89"),
  3723 => (x"d1",x"c4",x"91",x"bf"),
  3724 => (x"71",x"81",x"bf",x"cc"),
  3725 => (x"e4",x"d1",x"c4",x"1e"),
  3726 => (x"e0",x"c3",x"fd",x"49"),
  3727 => (x"c4",x"86",x"c4",x"87"),
  3728 => (x"c0",x"48",x"e8",x"f7"),
  3729 => (x"d1",x"f7",x"c4",x"78"),
  3730 => (x"c4",x"50",x"c1",x"48"),
  3731 => (x"c2",x"48",x"c4",x"f7"),
  3732 => (x"87",x"f9",x"cc",x"50"),
  3733 => (x"66",x"97",x"e4",x"c0"),
  3734 => (x"87",x"c9",x"c0",x"02"),
  3735 => (x"48",x"d0",x"f7",x"c4"),
  3736 => (x"e8",x"cc",x"50",x"c1"),
  3737 => (x"e8",x"49",x"c0",x"87"),
  3738 => (x"e0",x"cc",x"87",x"df"),
  3739 => (x"87",x"eb",x"ec",x"87"),
  3740 => (x"cc",x"02",x"98",x"70"),
  3741 => (x"e9",x"c0",x"87",x"d7"),
  3742 => (x"48",x"49",x"66",x"97"),
  3743 => (x"c0",x"98",x"c0",x"c3"),
  3744 => (x"70",x"58",x"a6",x"f0"),
  3745 => (x"dc",x"c0",x"02",x"98"),
  3746 => (x"c0",x"c1",x"48",x"87"),
  3747 => (x"a6",x"f0",x"c0",x"88"),
  3748 => (x"02",x"98",x"70",x"58"),
  3749 => (x"48",x"87",x"ed",x"c0"),
  3750 => (x"c0",x"88",x"c0",x"c1"),
  3751 => (x"70",x"58",x"a6",x"f0"),
  3752 => (x"cd",x"c1",x"02",x"98"),
  3753 => (x"97",x"e3",x"c0",x"87"),
  3754 => (x"31",x"d0",x"49",x"66"),
  3755 => (x"66",x"97",x"e4",x"c0"),
  3756 => (x"72",x"32",x"c8",x"4a"),
  3757 => (x"97",x"e5",x"c0",x"b1"),
  3758 => (x"71",x"48",x"4a",x"66"),
  3759 => (x"a6",x"f0",x"c0",x"b0"),
  3760 => (x"87",x"ff",x"c0",x"58"),
  3761 => (x"66",x"97",x"e4",x"c0"),
  3762 => (x"87",x"e7",x"e5",x"49"),
  3763 => (x"c0",x"1e",x"49",x"70"),
  3764 => (x"49",x"66",x"97",x"e7"),
  3765 => (x"70",x"87",x"dc",x"e5"),
  3766 => (x"ea",x"c0",x"1e",x"49"),
  3767 => (x"e5",x"49",x"66",x"97"),
  3768 => (x"4a",x"70",x"87",x"d1"),
  3769 => (x"c9",x"c4",x"ff",x"49"),
  3770 => (x"c0",x"86",x"c8",x"87"),
  3771 => (x"c0",x"58",x"a6",x"f0"),
  3772 => (x"e2",x"c0",x"87",x"d1"),
  3773 => (x"e5",x"49",x"66",x"97"),
  3774 => (x"ec",x"c0",x"87",x"d3"),
  3775 => (x"d1",x"c4",x"48",x"a6"),
  3776 => (x"c4",x"78",x"bf",x"d0"),
  3777 => (x"c0",x"48",x"c0",x"f7"),
  3778 => (x"d8",x"f7",x"c4",x"78"),
  3779 => (x"66",x"ec",x"c0",x"48"),
  3780 => (x"ed",x"e1",x"49",x"78"),
  3781 => (x"d8",x"f7",x"c4",x"87"),
  3782 => (x"ec",x"f7",x"c4",x"58"),
  3783 => (x"66",x"ec",x"c0",x"48"),
  3784 => (x"c0",x"d1",x"c4",x"40"),
  3785 => (x"f7",x"c4",x"78",x"bf"),
  3786 => (x"e1",x"c0",x"48",x"f8"),
  3787 => (x"c4",x"50",x"66",x"97"),
  3788 => (x"c1",x"48",x"f4",x"f7"),
  3789 => (x"f8",x"f7",x"c4",x"78"),
  3790 => (x"99",x"49",x"bf",x"97"),
  3791 => (x"87",x"c9",x"c0",x"05"),
  3792 => (x"48",x"c4",x"f7",x"c4"),
  3793 => (x"c6",x"c0",x"50",x"c4"),
  3794 => (x"c4",x"f7",x"c4",x"87"),
  3795 => (x"c0",x"50",x"c3",x"48"),
  3796 => (x"87",x"dc",x"e5",x"49"),
  3797 => (x"e9",x"87",x"f6",x"c8"),
  3798 => (x"98",x"70",x"87",x"c1"),
  3799 => (x"87",x"ed",x"c8",x"02"),
  3800 => (x"66",x"97",x"e9",x"c0"),
  3801 => (x"c0",x"c3",x"48",x"49"),
  3802 => (x"a6",x"f0",x"c0",x"98"),
  3803 => (x"02",x"98",x"70",x"58"),
  3804 => (x"48",x"87",x"dc",x"c0"),
  3805 => (x"c0",x"88",x"c0",x"c1"),
  3806 => (x"70",x"58",x"a6",x"f0"),
  3807 => (x"ed",x"c0",x"02",x"98"),
  3808 => (x"c0",x"c1",x"48",x"87"),
  3809 => (x"a6",x"f0",x"c0",x"88"),
  3810 => (x"02",x"98",x"70",x"58"),
  3811 => (x"c0",x"87",x"cd",x"c1"),
  3812 => (x"49",x"66",x"97",x"e3"),
  3813 => (x"e4",x"c0",x"31",x"d0"),
  3814 => (x"c8",x"4a",x"66",x"97"),
  3815 => (x"c0",x"b1",x"72",x"32"),
  3816 => (x"4a",x"66",x"97",x"e5"),
  3817 => (x"c0",x"b0",x"71",x"48"),
  3818 => (x"c1",x"58",x"a6",x"f0"),
  3819 => (x"e4",x"c0",x"87",x"f4"),
  3820 => (x"e1",x"49",x"66",x"97"),
  3821 => (x"49",x"70",x"87",x"fd"),
  3822 => (x"97",x"e7",x"c0",x"1e"),
  3823 => (x"f2",x"e1",x"49",x"66"),
  3824 => (x"1e",x"49",x"70",x"87"),
  3825 => (x"66",x"97",x"ea",x"c0"),
  3826 => (x"87",x"e7",x"e1",x"49"),
  3827 => (x"ff",x"49",x"4a",x"70"),
  3828 => (x"c8",x"87",x"df",x"c0"),
  3829 => (x"a6",x"f0",x"c0",x"86"),
  3830 => (x"87",x"c6",x"c1",x"58"),
  3831 => (x"66",x"97",x"e2",x"c0"),
  3832 => (x"87",x"cf",x"e1",x"49"),
  3833 => (x"c0",x"48",x"49",x"70"),
  3834 => (x"70",x"58",x"a6",x"f0"),
  3835 => (x"c6",x"c0",x"05",x"98"),
  3836 => (x"a6",x"ec",x"c0",x"87"),
  3837 => (x"c0",x"78",x"c1",x"48"),
  3838 => (x"c4",x"48",x"66",x"ec"),
  3839 => (x"b7",x"bf",x"c4",x"d1"),
  3840 => (x"cc",x"c0",x"06",x"a8"),
  3841 => (x"a6",x"f4",x"c0",x"87"),
  3842 => (x"c0",x"d1",x"c4",x"48"),
  3843 => (x"c9",x"c0",x"78",x"bf"),
  3844 => (x"a6",x"f4",x"c0",x"87"),
  3845 => (x"d4",x"d1",x"c4",x"48"),
  3846 => (x"ec",x"c0",x"78",x"bf"),
  3847 => (x"f4",x"c0",x"48",x"a6"),
  3848 => (x"f7",x"c4",x"78",x"66"),
  3849 => (x"e1",x"c0",x"48",x"f8"),
  3850 => (x"c4",x"50",x"66",x"97"),
  3851 => (x"c0",x"48",x"f0",x"f7"),
  3852 => (x"c4",x"78",x"66",x"ec"),
  3853 => (x"bf",x"97",x"f8",x"f7"),
  3854 => (x"c0",x"05",x"99",x"49"),
  3855 => (x"f7",x"c4",x"87",x"c9"),
  3856 => (x"50",x"c0",x"48",x"c4"),
  3857 => (x"c4",x"87",x"c6",x"c0"),
  3858 => (x"c3",x"48",x"c4",x"f7"),
  3859 => (x"f8",x"f7",x"c4",x"50"),
  3860 => (x"c2",x"49",x"bf",x"97"),
  3861 => (x"f4",x"c4",x"02",x"a9"),
  3862 => (x"e0",x"49",x"c0",x"87"),
  3863 => (x"ec",x"c4",x"87",x"eb"),
  3864 => (x"87",x"f7",x"e4",x"87"),
  3865 => (x"c4",x"02",x"98",x"70"),
  3866 => (x"f7",x"c4",x"87",x"e3"),
  3867 => (x"50",x"c4",x"48",x"c4"),
  3868 => (x"d4",x"e0",x"49",x"c0"),
  3869 => (x"87",x"d5",x"c4",x"87"),
  3870 => (x"70",x"87",x"e0",x"e4"),
  3871 => (x"cc",x"c4",x"02",x"98"),
  3872 => (x"d8",x"f7",x"c4",x"87"),
  3873 => (x"d1",x"c4",x"48",x"bf"),
  3874 => (x"c0",x"88",x"bf",x"d0"),
  3875 => (x"ca",x"58",x"a6",x"f0"),
  3876 => (x"a6",x"c1",x"7e",x"97"),
  3877 => (x"50",x"c0",x"c2",x"48"),
  3878 => (x"97",x"c4",x"f7",x"c4"),
  3879 => (x"f8",x"c0",x"48",x"bf"),
  3880 => (x"a8",x"c4",x"58",x"a6"),
  3881 => (x"87",x"c9",x"c0",x"05"),
  3882 => (x"48",x"a6",x"f4",x"c0"),
  3883 => (x"e1",x"c0",x"78",x"c2"),
  3884 => (x"66",x"f4",x"c0",x"87"),
  3885 => (x"05",x"a8",x"c3",x"48"),
  3886 => (x"c0",x"87",x"c9",x"c0"),
  3887 => (x"c0",x"48",x"a6",x"f8"),
  3888 => (x"87",x"c6",x"c0",x"78"),
  3889 => (x"48",x"a6",x"f8",x"c0"),
  3890 => (x"f4",x"c0",x"78",x"c3"),
  3891 => (x"f8",x"c0",x"48",x"a6"),
  3892 => (x"a6",x"c2",x"78",x"66"),
  3893 => (x"66",x"f4",x"c0",x"48"),
  3894 => (x"c4",x"50",x"c0",x"50"),
  3895 => (x"49",x"bf",x"d4",x"f7"),
  3896 => (x"dc",x"ff",x"81",x"c1"),
  3897 => (x"a6",x"c4",x"87",x"de"),
  3898 => (x"f7",x"c4",x"50",x"08"),
  3899 => (x"ff",x"49",x"bf",x"d4"),
  3900 => (x"c5",x"87",x"d1",x"dc"),
  3901 => (x"c0",x"50",x"08",x"a6"),
  3902 => (x"1e",x"4b",x"a6",x"f0"),
  3903 => (x"49",x"66",x"f0",x"c0"),
  3904 => (x"87",x"e4",x"fa",x"fe"),
  3905 => (x"66",x"97",x"f4",x"c0"),
  3906 => (x"f7",x"db",x"ff",x"49"),
  3907 => (x"08",x"a6",x"ca",x"87"),
  3908 => (x"97",x"f5",x"c0",x"50"),
  3909 => (x"db",x"ff",x"49",x"66"),
  3910 => (x"a6",x"cb",x"87",x"ea"),
  3911 => (x"f6",x"c0",x"50",x"08"),
  3912 => (x"ff",x"49",x"66",x"97"),
  3913 => (x"cc",x"87",x"dd",x"db"),
  3914 => (x"73",x"50",x"08",x"a6"),
  3915 => (x"d8",x"f7",x"c4",x"1e"),
  3916 => (x"f9",x"fe",x"49",x"bf"),
  3917 => (x"f8",x"c0",x"87",x"f2"),
  3918 => (x"ff",x"49",x"66",x"97"),
  3919 => (x"d1",x"87",x"c5",x"db"),
  3920 => (x"c0",x"50",x"08",x"a6"),
  3921 => (x"49",x"66",x"97",x"f9"),
  3922 => (x"87",x"f8",x"da",x"ff"),
  3923 => (x"50",x"08",x"a6",x"d2"),
  3924 => (x"66",x"97",x"fa",x"c0"),
  3925 => (x"eb",x"da",x"ff",x"49"),
  3926 => (x"08",x"a6",x"d3",x"87"),
  3927 => (x"ca",x"1e",x"c1",x"50"),
  3928 => (x"49",x"a6",x"d2",x"1e"),
  3929 => (x"87",x"d6",x"dd",x"ff"),
  3930 => (x"49",x"c0",x"86",x"d0"),
  3931 => (x"87",x"d9",x"dc",x"ff"),
  3932 => (x"c0",x"87",x"da",x"c0"),
  3933 => (x"e0",x"c0",x"1e",x"1e"),
  3934 => (x"ff",x"49",x"c5",x"1e"),
  3935 => (x"cc",x"87",x"f5",x"db"),
  3936 => (x"cc",x"f7",x"c4",x"86"),
  3937 => (x"c1",x"78",x"c0",x"48"),
  3938 => (x"fc",x"db",x"ff",x"49"),
  3939 => (x"8e",x"c4",x"ff",x"87"),
  3940 => (x"4c",x"26",x"4d",x"26"),
  3941 => (x"4f",x"26",x"4b",x"26"),
  3942 => (x"f4",x"1e",x"73",x"1e"),
  3943 => (x"4b",x"d4",x"ff",x"86"),
  3944 => (x"c8",x"48",x"d0",x"ff"),
  3945 => (x"e3",x"c1",x"78",x"c5"),
  3946 => (x"c0",x"4a",x"c0",x"7b"),
  3947 => (x"72",x"49",x"76",x"7b"),
  3948 => (x"c1",x"51",x"6b",x"81"),
  3949 => (x"aa",x"b7",x"ca",x"82"),
  3950 => (x"ff",x"87",x"f0",x"04"),
  3951 => (x"78",x"c4",x"48",x"d0"),
  3952 => (x"4b",x"26",x"8e",x"f4"),
  3953 => (x"c4",x"1e",x"4f",x"26"),
  3954 => (x"c1",x"48",x"d1",x"f7"),
  3955 => (x"1e",x"4f",x"26",x"50"),
  3956 => (x"48",x"c0",x"f7",x"c4"),
  3957 => (x"f7",x"c4",x"78",x"c0"),
  3958 => (x"40",x"c0",x"48",x"d4"),
  3959 => (x"e0",x"f7",x"c4",x"78"),
  3960 => (x"c4",x"78",x"c0",x"48"),
  3961 => (x"c1",x"48",x"c5",x"f7"),
  3962 => (x"ec",x"d1",x"c4",x"50"),
  3963 => (x"87",x"c4",x"02",x"bf"),
  3964 => (x"87",x"c2",x"49",x"c0"),
  3965 => (x"f7",x"c4",x"49",x"c1"),
  3966 => (x"c4",x"59",x"97",x"c8"),
  3967 => (x"c0",x"48",x"e4",x"f7"),
  3968 => (x"f7",x"c4",x"78",x"40"),
  3969 => (x"40",x"c0",x"48",x"cc"),
  3970 => (x"f7",x"c4",x"50",x"50"),
  3971 => (x"40",x"c0",x"48",x"ec"),
  3972 => (x"f8",x"f7",x"c4",x"78"),
  3973 => (x"c4",x"50",x"c0",x"48"),
  3974 => (x"c0",x"48",x"fa",x"f7"),
  3975 => (x"f7",x"c4",x"78",x"9f"),
  3976 => (x"50",x"c1",x"48",x"d2"),
  3977 => (x"73",x"1e",x"4f",x"26"),
  3978 => (x"48",x"d0",x"ff",x"1e"),
  3979 => (x"ff",x"78",x"c5",x"c8"),
  3980 => (x"e0",x"c1",x"48",x"d4"),
  3981 => (x"c3",x"49",x"68",x"78"),
  3982 => (x"d0",x"ff",x"99",x"ff"),
  3983 => (x"71",x"78",x"c4",x"48"),
  3984 => (x"99",x"c1",x"49",x"4b"),
  3985 => (x"e6",x"87",x"c3",x"02"),
  3986 => (x"49",x"73",x"87",x"c0"),
  3987 => (x"c3",x"02",x"99",x"c2"),
  3988 => (x"87",x"c4",x"fd",x"87"),
  3989 => (x"99",x"c4",x"49",x"73"),
  3990 => (x"fd",x"87",x"c3",x"02"),
  3991 => (x"49",x"73",x"87",x"e8"),
  3992 => (x"d6",x"02",x"99",x"c8"),
  3993 => (x"87",x"e7",x"fd",x"87"),
  3994 => (x"c8",x"48",x"d0",x"ff"),
  3995 => (x"d4",x"ff",x"78",x"c5"),
  3996 => (x"78",x"e6",x"c1",x"48"),
  3997 => (x"d0",x"ff",x"78",x"c0"),
  3998 => (x"73",x"78",x"c4",x"48"),
  3999 => (x"c4",x"99",x"d0",x"49"),
  4000 => (x"59",x"97",x"d6",x"f7"),
  4001 => (x"87",x"fa",x"dc",x"ff"),
  4002 => (x"bf",x"cc",x"f7",x"c4"),
  4003 => (x"c4",x"87",x"d7",x"02"),
  4004 => (x"05",x"bf",x"c0",x"f7"),
  4005 => (x"f7",x"c4",x"87",x"d0"),
  4006 => (x"49",x"bf",x"9f",x"fa"),
  4007 => (x"87",x"e9",x"d7",x"ff"),
  4008 => (x"48",x"cc",x"f7",x"c4"),
  4009 => (x"f7",x"c4",x"78",x"c0"),
  4010 => (x"02",x"bf",x"97",x"d0"),
  4011 => (x"d0",x"ff",x"87",x"d9"),
  4012 => (x"78",x"c5",x"c8",x"48"),
  4013 => (x"c1",x"48",x"d4",x"ff"),
  4014 => (x"78",x"c0",x"78",x"e5"),
  4015 => (x"c4",x"48",x"d0",x"ff"),
  4016 => (x"d0",x"f7",x"c4",x"78"),
  4017 => (x"26",x"50",x"c0",x"48"),
  4018 => (x"00",x"4f",x"26",x"4b"),
  4019 => (x"00",x"00",x"00",x"00"),
  4020 => (x"ff",x"4a",x"71",x"1e"),
  4021 => (x"72",x"49",x"bf",x"c8"),
  4022 => (x"4f",x"26",x"48",x"a1"),
  4023 => (x"bf",x"c8",x"ff",x"1e"),
  4024 => (x"c0",x"c0",x"fe",x"89"),
  4025 => (x"a9",x"c0",x"c0",x"c0"),
  4026 => (x"c0",x"87",x"c4",x"01"),
  4027 => (x"c1",x"87",x"c2",x"4a"),
  4028 => (x"26",x"48",x"72",x"4a"),
  4029 => (x"fd",x"c3",x"1e",x"4f"),
  4030 => (x"c1",x"49",x"bf",x"c4"),
  4031 => (x"c8",x"fd",x"c3",x"b9"),
  4032 => (x"48",x"d4",x"ff",x"59"),
  4033 => (x"ff",x"78",x"ff",x"c3"),
  4034 => (x"e1",x"c0",x"48",x"d0"),
  4035 => (x"48",x"d4",x"ff",x"78"),
  4036 => (x"31",x"c4",x"78",x"c1"),
  4037 => (x"d0",x"ff",x"78",x"71"),
  4038 => (x"78",x"e0",x"c0",x"48"),
  4039 => (x"c3",x"1e",x"4f",x"26"),
  4040 => (x"c4",x"1e",x"f8",x"fc"),
  4041 => (x"fc",x"49",x"e8",x"cb"),
  4042 => (x"c4",x"87",x"dc",x"e9"),
  4043 => (x"02",x"98",x"70",x"86"),
  4044 => (x"c0",x"ff",x"87",x"c3"),
  4045 => (x"00",x"4f",x"26",x"87"),
  4046 => (x"48",x"4b",x"35",x"31"),
  4047 => (x"20",x"20",x"20",x"5a"),
  4048 => (x"00",x"47",x"46",x"43"),
  4049 => (x"00",x"00",x"00",x"00"),
  4050 => (x"dc",x"f2",x"c1",x"1e"),
  4051 => (x"c1",x"50",x"c1",x"48"),
  4052 => (x"c1",x"48",x"cc",x"c6"),
  4053 => (x"f4",x"fd",x"c3",x"50"),
  4054 => (x"c8",x"fd",x"49",x"bf"),
  4055 => (x"48",x"c0",x"87",x"ef"),
  4056 => (x"00",x"00",x"4f",x"26"),
  4057 => (x"11",x"14",x"12",x"58"),
  4058 => (x"23",x"1c",x"1b",x"1d"),
  4059 => (x"91",x"94",x"59",x"5a"),
  4060 => (x"f4",x"eb",x"f2",x"f5"),
  4061 => (x"00",x"00",x"3f",x"78"),
  4062 => (x"4f",x"54",x"55",x"41"),
  4063 => (x"54",x"4f",x"4f",x"42"),
  4064 => (x"00",x"58",x"47",x"53"),
		others => (others => x"00")
	);
	signal q1_local : word_t;

	-- Altera Quartus attributes
	attribute ramstyle: string;
	attribute ramstyle of ram: signal is "no_rw_check";

begin  -- rtl

	addr1 <= to_integer(unsigned(addr(ADDR_WIDTH-1 downto 0)));

	-- Reorganize the read data from the RAM to match the output
	q(7 downto 0) <= q1_local(3);
	q(15 downto 8) <= q1_local(2);
	q(23 downto 16) <= q1_local(1);
	q(31 downto 24) <= q1_local(0);

	process(clk)
	begin
		if(rising_edge(clk)) then 
			if(we = '1') then
				-- edit this code if using other than four bytes per word
				if (bytesel(3) = '1') then
					ram(addr1)(3) <= d(7 downto 0);
				end if;
				if (bytesel(2) = '1') then
					ram(addr1)(2) <= d(15 downto 8);
				end if;
				if (bytesel(1) = '1') then
					ram(addr1)(1) <= d(23 downto 16);
				end if;
				if (bytesel(0) = '1') then
					ram(addr1)(0) <= d(31 downto 24);
				end if;
			end if;
			q1_local <= ram(addr1);
		end if;
	end process;
  
end rtl;

