library ieee;
use ieee.std_logic_1164.all;
use ieee.numeric_std.all;

entity controller_rom1 is
generic	(
	ADDR_WIDTH : integer := 8; -- ROM's address width (words, not bytes)
	COL_WIDTH  : integer := 8;  -- Column width (8bit -> byte)
	NB_COL     : integer := 4  -- Number of columns in memory
	);
port (
	clk : in std_logic;
	reset_n : in std_logic := '1';
	addr : in std_logic_vector(ADDR_WIDTH-1 downto 0);
	q : out std_logic_vector(31 downto 0);
	-- Allow writes - defaults supplied to simplify projects that don't need to write.
	d : in std_logic_vector(31 downto 0) := X"00000000";
	we : in std_logic := '0';
	bytesel : in std_logic_vector(3 downto 0) := "1111"
);
end entity;

architecture arch of controller_rom1 is

-- type word_t is std_logic_vector(31 downto 0);
type ram_type is array (0 to 2 ** ADDR_WIDTH - 1) of std_logic_vector(NB_COL * COL_WIDTH - 1 downto 0);

signal ram : ram_type :=
(

     0 => x"0487da01",
     1 => x"580e87dd",
     2 => x"0e5a595e",
     3 => x"00002927",
     4 => x"4a260f00",
     5 => x"48264926",
     6 => x"082680ff",
     7 => x"002d274f",
     8 => x"274f0000",
     9 => x"0000002a",
    10 => x"fd004f4f",
    11 => x"fcf7c487",
    12 => x"86c0c54e",
    13 => x"49fcf7c4",
    14 => x"48c4fec3",
    15 => x"4040c089",
    16 => x"89d04040",
    17 => x"c187f603",
    18 => x"0087faf0",
    19 => x"1e87fc98",
    20 => x"48121e72",
    21 => x"87c40211",
    22 => x"87f60288",
    23 => x"4f264a26",
    24 => x"731e721e",
    25 => x"1148121e",
    26 => x"4b87ca02",
    27 => x"9b98dfc3",
    28 => x"f0028873",
    29 => x"264b2687",
    30 => x"1e4f264a",
    31 => x"1e721e73",
    32 => x"ca048bc1",
    33 => x"11481287",
    34 => x"8887c402",
    35 => x"2687f102",
    36 => x"264b264a",
    37 => x"1e741e4f",
    38 => x"1e721e73",
    39 => x"d0048bc1",
    40 => x"11481287",
    41 => x"4c87ca02",
    42 => x"9c98dfc3",
    43 => x"eb028874",
    44 => x"264a2687",
    45 => x"264c264b",
    46 => x"48731e4f",
    47 => x"02a97381",
    48 => x"531287c5",
    49 => x"2687f605",
    50 => x"48731e4f",
    51 => x"05a97381",
    52 => x"87f95372",
    53 => x"5e0e4f26",
    54 => x"0e5d5c5b",
    55 => x"4d7186f4",
    56 => x"c048a6c4",
    57 => x"4b66dc78",
    58 => x"c048a6c8",
    59 => x"7e971578",
    60 => x"c0026e97",
    61 => x"4c1387f0",
    62 => x"87da029c",
    63 => x"744a6e97",
    64 => x"05aab749",
    65 => x"a6c887c9",
    66 => x"c078c148",
    67 => x"1387c24c",
    68 => x"059c744c",
    69 => x"66c887e6",
    70 => x"c487cb02",
    71 => x"80c14866",
    72 => x"fe58a6c8",
    73 => x"66c487ff",
    74 => x"268ef448",
    75 => x"264c264d",
    76 => x"1e4f264b",
    77 => x"c1c14a71",
    78 => x"d904aab7",
    79 => x"b7c6c187",
    80 => x"87d201aa",
    81 => x"d04866c4",
    82 => x"87ca05a8",
    83 => x"f7c04972",
    84 => x"c0487189",
    85 => x"e1c187ec",
    86 => x"d804aab7",
    87 => x"b7e6c187",
    88 => x"87d101aa",
    89 => x"d04866c4",
    90 => x"87c905a8",
    91 => x"d7c14972",
    92 => x"cd487189",
    93 => x"8af0c087",
    94 => x"06aab7c9",
    95 => x"4aff87c2",
    96 => x"4f264872",
    97 => x"5c5b5e0e",
    98 => x"86f80e5d",
    99 => x"a6c47e71",
   100 => x"4c78c048",
   101 => x"1ea7f9c1",
   102 => x"fc4966c4",
   103 => x"86c487f8",
   104 => x"4b6e4970",
   105 => x"6b978371",
   106 => x"a9edc049",
   107 => x"c487c605",
   108 => x"78c148a6",
   109 => x"0266d883",
   110 => x"66d887c5",
   111 => x"970b7b0b",
   112 => x"87d3056b",
   113 => x"c70266c4",
   114 => x"c04a7487",
   115 => x"87c28a0a",
   116 => x"48724a74",
   117 => x"dc87efc0",
   118 => x"49131e66",
   119 => x"c487d4fd",
   120 => x"c04d7086",
   121 => x"d403adb7",
   122 => x"0266c487",
   123 => x"487487c9",
   124 => x"708808c0",
   125 => x"7487c27e",
   126 => x"c9486e7e",
   127 => x"9466dc87",
   128 => x"fe4ca475",
   129 => x"8ef887ef",
   130 => x"4c264d26",
   131 => x"4f264b26",
   132 => x"731e0020",
   133 => x"029a721e",
   134 => x"c087e7c0",
   135 => x"724bc148",
   136 => x"87d106a9",
   137 => x"c9068272",
   138 => x"72837387",
   139 => x"87f401a9",
   140 => x"b2c187c3",
   141 => x"03a9723a",
   142 => x"07807389",
   143 => x"052b2ac1",
   144 => x"4b2687f3",
   145 => x"751e4f26",
   146 => x"714dc41e",
   147 => x"ff04a1b7",
   148 => x"c381c1b9",
   149 => x"b77207bd",
   150 => x"baff04a2",
   151 => x"bdc182c1",
   152 => x"87eefe07",
   153 => x"ff042dc1",
   154 => x"0780c1b8",
   155 => x"b9ff042d",
   156 => x"260781c1",
   157 => x"1e4f264d",
   158 => x"4a711e73",
   159 => x"494b66c8",
   160 => x"99718bc1",
   161 => x"1287cf02",
   162 => x"08d4ff48",
   163 => x"c1497378",
   164 => x"0599718b",
   165 => x"4b2687f1",
   166 => x"5e0e4f26",
   167 => x"710e5c5b",
   168 => x"4cd4ff4a",
   169 => x"494b66cc",
   170 => x"99718bc1",
   171 => x"c387ce02",
   172 => x"526c7cff",
   173 => x"8bc14973",
   174 => x"f2059971",
   175 => x"264c2687",
   176 => x"1e4f264b",
   177 => x"d4ff1e73",
   178 => x"7bffc34b",
   179 => x"ffc34a6b",
   180 => x"c8496b7b",
   181 => x"c3b17232",
   182 => x"4a6b7bff",
   183 => x"b27131c8",
   184 => x"6b7bffc3",
   185 => x"7232c849",
   186 => x"264871b1",
   187 => x"0e4f264b",
   188 => x"5d5c5b5e",
   189 => x"ff4d710e",
   190 => x"49754cd4",
   191 => x"7199ffc3",
   192 => x"c4fec37c",
   193 => x"87c805bf",
   194 => x"c94866d0",
   195 => x"58a6d430",
   196 => x"d84966d0",
   197 => x"99ffc329",
   198 => x"66d07c71",
   199 => x"c329d049",
   200 => x"7c7199ff",
   201 => x"c84966d0",
   202 => x"99ffc329",
   203 => x"66d07c71",
   204 => x"99ffc349",
   205 => x"49757c71",
   206 => x"ffc329d0",
   207 => x"6c7c7199",
   208 => x"fff0c94b",
   209 => x"abffc34a",
   210 => x"4987cf05",
   211 => x"4b6c7c71",
   212 => x"c5028ac1",
   213 => x"02ab7187",
   214 => x"487387f2",
   215 => x"4c264d26",
   216 => x"4f264b26",
   217 => x"ff49c01e",
   218 => x"ffc348d4",
   219 => x"c381c178",
   220 => x"04a9b7c8",
   221 => x"4f2687f1",
   222 => x"5c5b5e0e",
   223 => x"ffc00e5d",
   224 => x"4df7c1f0",
   225 => x"c0c0c0c1",
   226 => x"ff4bc0c0",
   227 => x"f8c487d6",
   228 => x"1ec04cdf",
   229 => x"d6fd4975",
   230 => x"c186c487",
   231 => x"e5c005a8",
   232 => x"48d4ff87",
   233 => x"7378ffc3",
   234 => x"f0e1c01e",
   235 => x"fc49e9c1",
   236 => x"86c487fd",
   237 => x"ca059870",
   238 => x"48d4ff87",
   239 => x"c178ffc3",
   240 => x"fe87cb48",
   241 => x"8cc187de",
   242 => x"87c6ff05",
   243 => x"4d2648c0",
   244 => x"4b264c26",
   245 => x"5e0e4f26",
   246 => x"c00e5c5b",
   247 => x"c1c1f0ff",
   248 => x"48d4ff4c",
   249 => x"d378ffc3",
   250 => x"741ec04b",
   251 => x"87fffb49",
   252 => x"987086c4",
   253 => x"ff87ca05",
   254 => x"ffc348d4",
   255 => x"ca48c178",
   256 => x"87e0fd87",
   257 => x"e0058bc1",
   258 => x"2648c087",
   259 => x"264b264c",
   260 => x"5b5e0e4f",
   261 => x"c30e5d5c",
   262 => x"d4ff4dff",
   263 => x"87c4fd4b",
   264 => x"c01eeac6",
   265 => x"c8c1f0e1",
   266 => x"87c3fb49",
   267 => x"a8c186c4",
   268 => x"fe87c802",
   269 => x"48c087e0",
   270 => x"fa87e2c1",
   271 => x"497087c5",
   272 => x"99ffffcf",
   273 => x"02a9eac6",
   274 => x"c9fe87c8",
   275 => x"c148c087",
   276 => x"7b7587cb",
   277 => x"fc4cf1c0",
   278 => x"987087de",
   279 => x"87ecc002",
   280 => x"ffc01ec0",
   281 => x"49fac1f0",
   282 => x"c487c4fa",
   283 => x"05987086",
   284 => x"7b7587da",
   285 => x"7b75496b",
   286 => x"7b757b75",
   287 => x"c0c17b75",
   288 => x"87c40299",
   289 => x"87d548c1",
   290 => x"87d148c0",
   291 => x"c405acc2",
   292 => x"c848c087",
   293 => x"058cc187",
   294 => x"c087fcfe",
   295 => x"264d2648",
   296 => x"264b264c",
   297 => x"5b5e0e4f",
   298 => x"ff0e5d5c",
   299 => x"e5c04dd0",
   300 => x"4cc0c1d0",
   301 => x"48c4fec3",
   302 => x"4bc778c1",
   303 => x"e3fa7dc2",
   304 => x"c07dc387",
   305 => x"f849741e",
   306 => x"86c487e5",
   307 => x"c105a8c1",
   308 => x"abc24b87",
   309 => x"c087c505",
   310 => x"87f6c048",
   311 => x"ff058bc1",
   312 => x"ecfc87da",
   313 => x"c8fec387",
   314 => x"05987058",
   315 => x"1ec187cd",
   316 => x"c1f0ffc0",
   317 => x"f6f749d0",
   318 => x"ff86c487",
   319 => x"ffc348d4",
   320 => x"87c3c378",
   321 => x"58ccfec3",
   322 => x"d4ff7dc2",
   323 => x"78ffc348",
   324 => x"4d2648c1",
   325 => x"4b264c26",
   326 => x"5e0e4f26",
   327 => x"0e5d5c5b",
   328 => x"4b7186fc",
   329 => x"c04cd4ff",
   330 => x"cdeec57e",
   331 => x"ffc34adf",
   332 => x"c3496c7c",
   333 => x"c005a9fe",
   334 => x"4d7487f8",
   335 => x"cc029b73",
   336 => x"1e66d487",
   337 => x"d1f54973",
   338 => x"d486c487",
   339 => x"48d0ff87",
   340 => x"d478d1c4",
   341 => x"ffc34a66",
   342 => x"058ac17d",
   343 => x"a6d887f8",
   344 => x"7cffc35a",
   345 => x"059b737c",
   346 => x"d0ff87c5",
   347 => x"c178d048",
   348 => x"8ac17e4a",
   349 => x"87f6fe05",
   350 => x"8efc486e",
   351 => x"4c264d26",
   352 => x"4f264b26",
   353 => x"711e731e",
   354 => x"ff4bc04a",
   355 => x"ffc348d4",
   356 => x"48d0ff78",
   357 => x"ff78c3c4",
   358 => x"ffc348d4",
   359 => x"c01e7278",
   360 => x"d1c1f0ff",
   361 => x"87c7f549",
   362 => x"987086c4",
   363 => x"c887d205",
   364 => x"66cc1ec0",
   365 => x"87e2fd49",
   366 => x"4b7086c4",
   367 => x"c248d0ff",
   368 => x"26487378",
   369 => x"0e4f264b",
   370 => x"5d5c5b5e",
   371 => x"c01ec00e",
   372 => x"c9c1f0ff",
   373 => x"87d7f449",
   374 => x"fec31ed2",
   375 => x"f9fc49cc",
   376 => x"c086c887",
   377 => x"d284c14c",
   378 => x"f804acb7",
   379 => x"ccfec387",
   380 => x"c349bf97",
   381 => x"c0c199c0",
   382 => x"e7c005a9",
   383 => x"d3fec387",
   384 => x"d049bf97",
   385 => x"d4fec331",
   386 => x"c84abf97",
   387 => x"c3b17232",
   388 => x"bf97d5fe",
   389 => x"4c71b14a",
   390 => x"ffffffcf",
   391 => x"ca84c19c",
   392 => x"87e7c134",
   393 => x"97d5fec3",
   394 => x"31c149bf",
   395 => x"fec399c6",
   396 => x"4abf97d6",
   397 => x"722ab7c7",
   398 => x"d1fec3b1",
   399 => x"4d4abf97",
   400 => x"fec39dcf",
   401 => x"4abf97d2",
   402 => x"32ca9ac3",
   403 => x"97d3fec3",
   404 => x"33c24bbf",
   405 => x"fec3b273",
   406 => x"4bbf97d4",
   407 => x"c69bc0c3",
   408 => x"b2732bb7",
   409 => x"48c181c2",
   410 => x"49703071",
   411 => x"307548c1",
   412 => x"4c724d70",
   413 => x"947184c1",
   414 => x"adb7c0c8",
   415 => x"c187cc06",
   416 => x"c82db734",
   417 => x"01adb7c0",
   418 => x"7487f4ff",
   419 => x"264d2648",
   420 => x"264b264c",
   421 => x"5b5e0e4f",
   422 => x"f80e5d5c",
   423 => x"f4c6c486",
   424 => x"c378c048",
   425 => x"c01eecfe",
   426 => x"87d8fb49",
   427 => x"987086c4",
   428 => x"c087c505",
   429 => x"87cec948",
   430 => x"7ec14dc0",
   431 => x"bfe0fec0",
   432 => x"e2ffc349",
   433 => x"4bc8714a",
   434 => x"7087f0e6",
   435 => x"87c20598",
   436 => x"fec07ec0",
   437 => x"c349bfdc",
   438 => x"714afeff",
   439 => x"dae64bc8",
   440 => x"05987087",
   441 => x"7ec087c2",
   442 => x"fdc0026e",
   443 => x"f2c5c487",
   444 => x"c6c44dbf",
   445 => x"7ebf9fea",
   446 => x"ead6c548",
   447 => x"87c705a8",
   448 => x"bff2c5c4",
   449 => x"6e87ce4d",
   450 => x"d5e9ca48",
   451 => x"87c502a8",
   452 => x"f1c748c0",
   453 => x"ecfec387",
   454 => x"f949751e",
   455 => x"86c487e6",
   456 => x"c5059870",
   457 => x"c748c087",
   458 => x"fec087dc",
   459 => x"c349bfdc",
   460 => x"714afeff",
   461 => x"c2e54bc8",
   462 => x"05987087",
   463 => x"c6c487c8",
   464 => x"78c148f4",
   465 => x"fec087da",
   466 => x"c349bfe0",
   467 => x"714ae2ff",
   468 => x"e6e44bc8",
   469 => x"02987087",
   470 => x"c087c5c0",
   471 => x"87e6c648",
   472 => x"97eac6c4",
   473 => x"d5c149bf",
   474 => x"cdc005a9",
   475 => x"ebc6c487",
   476 => x"c249bf97",
   477 => x"c002a9ea",
   478 => x"48c087c5",
   479 => x"c387c7c6",
   480 => x"bf97ecfe",
   481 => x"e9c3487e",
   482 => x"cec002a8",
   483 => x"c3486e87",
   484 => x"c002a8eb",
   485 => x"48c087c5",
   486 => x"c387ebc5",
   487 => x"bf97f7fe",
   488 => x"c0059949",
   489 => x"fec387cc",
   490 => x"49bf97f8",
   491 => x"c002a9c2",
   492 => x"48c087c5",
   493 => x"c387cfc5",
   494 => x"bf97f9fe",
   495 => x"f0c6c448",
   496 => x"484c7058",
   497 => x"c6c488c1",
   498 => x"fec358f4",
   499 => x"49bf97fa",
   500 => x"fec38175",
   501 => x"4abf97fb",
   502 => x"a17232c8",
   503 => x"c4cbc47e",
   504 => x"c3786e48",
   505 => x"bf97fcfe",
   506 => x"58a6c848",
   507 => x"bff4c6c4",
   508 => x"87d4c202",
   509 => x"bfdcfec0",
   510 => x"feffc349",
   511 => x"4bc8714a",
   512 => x"7087f8e1",
   513 => x"c5c00298",
   514 => x"c348c087",
   515 => x"c6c487f8",
   516 => x"c44cbfec",
   517 => x"c35cd8cb",
   518 => x"bf97d1ff",
   519 => x"c331c849",
   520 => x"bf97d0ff",
   521 => x"c349a14a",
   522 => x"bf97d2ff",
   523 => x"7232d04a",
   524 => x"ffc349a1",
   525 => x"4abf97d3",
   526 => x"a17232d8",
   527 => x"9166c449",
   528 => x"bfc4cbc4",
   529 => x"cccbc481",
   530 => x"d9ffc359",
   531 => x"c84abf97",
   532 => x"d8ffc332",
   533 => x"a24bbf97",
   534 => x"daffc34a",
   535 => x"d04bbf97",
   536 => x"4aa27333",
   537 => x"97dbffc3",
   538 => x"9bcf4bbf",
   539 => x"a27333d8",
   540 => x"d0cbc44a",
   541 => x"cccbc45a",
   542 => x"8ac24abf",
   543 => x"cbc49274",
   544 => x"a17248d0",
   545 => x"87cac178",
   546 => x"97fefec3",
   547 => x"31c849bf",
   548 => x"97fdfec3",
   549 => x"49a14abf",
   550 => x"59fcc6c4",
   551 => x"bff8c6c4",
   552 => x"c731c549",
   553 => x"29c981ff",
   554 => x"59d8cbc4",
   555 => x"97c3ffc3",
   556 => x"32c84abf",
   557 => x"97c2ffc3",
   558 => x"4aa24bbf",
   559 => x"6e9266c4",
   560 => x"d4cbc482",
   561 => x"cccbc45a",
   562 => x"c478c048",
   563 => x"7248c8cb",
   564 => x"cbc478a1",
   565 => x"cbc448d8",
   566 => x"c478bfcc",
   567 => x"c448dccb",
   568 => x"78bfd0cb",
   569 => x"bff4c6c4",
   570 => x"87c9c002",
   571 => x"30c44874",
   572 => x"c9c07e70",
   573 => x"d4cbc487",
   574 => x"30c448bf",
   575 => x"c6c47e70",
   576 => x"786e48f8",
   577 => x"8ef848c1",
   578 => x"4c264d26",
   579 => x"4f264b26",
   580 => x"5c5b5e0e",
   581 => x"4a710e5d",
   582 => x"bff4c6c4",
   583 => x"7287cb02",
   584 => x"722bc74b",
   585 => x"9cffc14c",
   586 => x"4b7287c9",
   587 => x"4c722bc8",
   588 => x"c49cffc3",
   589 => x"83bfc4cb",
   590 => x"bfd8fec0",
   591 => x"87d902ab",
   592 => x"5bdcfec0",
   593 => x"1eecfec3",
   594 => x"f7f04973",
   595 => x"7086c487",
   596 => x"87c50598",
   597 => x"e6c048c0",
   598 => x"f4c6c487",
   599 => x"87d202bf",
   600 => x"91c44974",
   601 => x"81ecfec3",
   602 => x"ffcf4d69",
   603 => x"9dffffff",
   604 => x"497487cb",
   605 => x"fec391c2",
   606 => x"699f81ec",
   607 => x"2648754d",
   608 => x"264c264d",
   609 => x"0e4f264b",
   610 => x"5d5c5b5e",
   611 => x"cc86f40e",
   612 => x"66c859a6",
   613 => x"c087c505",
   614 => x"87c8c348",
   615 => x"c84866c8",
   616 => x"6e7e7080",
   617 => x"dc78c048",
   618 => x"87c70266",
   619 => x"bf9766dc",
   620 => x"c087c505",
   621 => x"87ecc248",
   622 => x"49c11ec0",
   623 => x"c487dbcf",
   624 => x"9c4c7086",
   625 => x"87fcc002",
   626 => x"4afcc6c4",
   627 => x"ff4966dc",
   628 => x"7087cdda",
   629 => x"ebc00298",
   630 => x"dc4a7487",
   631 => x"4bcb4966",
   632 => x"87f1daff",
   633 => x"db029870",
   634 => x"741ec087",
   635 => x"87c4029c",
   636 => x"87c24dc0",
   637 => x"49754dc1",
   638 => x"c487dfce",
   639 => x"9c4c7086",
   640 => x"87c4ff05",
   641 => x"c1029c74",
   642 => x"a4dc87d8",
   643 => x"69486e49",
   644 => x"49a4da78",
   645 => x"c44866c8",
   646 => x"58a6c880",
   647 => x"c448699f",
   648 => x"c4780866",
   649 => x"02bff4c6",
   650 => x"a4d487d2",
   651 => x"49699f49",
   652 => x"99ffffc0",
   653 => x"30d04871",
   654 => x"87c27e70",
   655 => x"496e7ec0",
   656 => x"bf66c448",
   657 => x"0866c480",
   658 => x"4866c878",
   659 => x"66c878c0",
   660 => x"c481cc49",
   661 => x"c879bf66",
   662 => x"81d04966",
   663 => x"48c179c0",
   664 => x"48c087c2",
   665 => x"4d268ef4",
   666 => x"4b264c26",
   667 => x"5e0e4f26",
   668 => x"0e5d5c5b",
   669 => x"029c4c71",
   670 => x"c887cac1",
   671 => x"026949a4",
   672 => x"d087c2c1",
   673 => x"496c4a66",
   674 => x"5aa6d482",
   675 => x"b94d66d0",
   676 => x"bff0c6c4",
   677 => x"72baff4a",
   678 => x"02997199",
   679 => x"c487e4c0",
   680 => x"496b4ba4",
   681 => x"7087e9f9",
   682 => x"ecc6c47b",
   683 => x"816c49bf",
   684 => x"b9757c71",
   685 => x"bff0c6c4",
   686 => x"72baff4a",
   687 => x"05997199",
   688 => x"7587dcff",
   689 => x"264d267c",
   690 => x"264b264c",
   691 => x"1e731e4f",
   692 => x"029b4b71",
   693 => x"a3c887c7",
   694 => x"c5056949",
   695 => x"c048c087",
   696 => x"cbc487f7",
   697 => x"c44abfc8",
   698 => x"496949a3",
   699 => x"c6c489c2",
   700 => x"7191bfec",
   701 => x"c6c44aa2",
   702 => x"6b49bff0",
   703 => x"4aa27199",
   704 => x"5adcfec0",
   705 => x"721e66c8",
   706 => x"87f8e949",
   707 => x"987086c4",
   708 => x"c087c405",
   709 => x"c187c248",
   710 => x"264b2648",
   711 => x"5b5e0e4f",
   712 => x"fc0e5d5c",
   713 => x"d44b7186",
   714 => x"9b734d66",
   715 => x"87ccc102",
   716 => x"6949a3c8",
   717 => x"87c4c102",
   718 => x"c44ca3d0",
   719 => x"49bff0c6",
   720 => x"4a6cb9ff",
   721 => x"66d47e99",
   722 => x"87cd06a9",
   723 => x"cc7c7bc0",
   724 => x"a3c44aa3",
   725 => x"ca796a49",
   726 => x"f8497287",
   727 => x"66d499c0",
   728 => x"758d714d",
   729 => x"7129c949",
   730 => x"fc49731e",
   731 => x"fec387c0",
   732 => x"49731eec",
   733 => x"c887d6fd",
   734 => x"7c66d486",
   735 => x"4d268efc",
   736 => x"4b264c26",
   737 => x"5e0e4f26",
   738 => x"0e5d5c5b",
   739 => x"a6d086f0",
   740 => x"66e0c059",
   741 => x"66e4c04c",
   742 => x"0266cc4b",
   743 => x"c84887ca",
   744 => x"6e7e7080",
   745 => x"87c505bf",
   746 => x"ecc348c0",
   747 => x"4d66cc87",
   748 => x"497385d0",
   749 => x"6d48a6c4",
   750 => x"8166c478",
   751 => x"bf6e80c4",
   752 => x"a966c878",
   753 => x"4987c606",
   754 => x"718966c4",
   755 => x"abb7c04b",
   756 => x"4887c401",
   757 => x"c487c2c3",
   758 => x"ffc74866",
   759 => x"6e7e7098",
   760 => x"87cdc102",
   761 => x"6e49c0c8",
   762 => x"59a6cc89",
   763 => x"4aecfec3",
   764 => x"66c8826e",
   765 => x"c303abb7",
   766 => x"5ba6cc87",
   767 => x"484966c8",
   768 => x"708066c4",
   769 => x"8b66c87d",
   770 => x"88c14849",
   771 => x"7158a6cc",
   772 => x"87d30299",
   773 => x"c17c9712",
   774 => x"4966c884",
   775 => x"cc88c148",
   776 => x"997158a6",
   777 => x"c187ed05",
   778 => x"4966d01e",
   779 => x"c487fff8",
   780 => x"abb7c086",
   781 => x"87dfc106",
   782 => x"abb7ffc7",
   783 => x"87e2c006",
   784 => x"66d01e74",
   785 => x"87c5fa49",
   786 => x"6d84c0c8",
   787 => x"80c0c848",
   788 => x"c0c87d70",
   789 => x"d41ec18b",
   790 => x"d1f84966",
   791 => x"c086c887",
   792 => x"fec387ee",
   793 => x"66d01eec",
   794 => x"87e1f949",
   795 => x"fec386c4",
   796 => x"49734aec",
   797 => x"70806d48",
   798 => x"c149737d",
   799 => x"0299718b",
   800 => x"971287ce",
   801 => x"7384c17c",
   802 => x"718bc149",
   803 => x"87f20599",
   804 => x"01abb7c0",
   805 => x"c187e1fe",
   806 => x"268ef048",
   807 => x"264c264d",
   808 => x"0e4f264b",
   809 => x"5d5c5b5e",
   810 => x"9b4b710e",
   811 => x"c887c702",
   812 => x"056d4da3",
   813 => x"48ff87c5",
   814 => x"d087fdc0",
   815 => x"496c4ca3",
   816 => x"0599ffc7",
   817 => x"026c87d8",
   818 => x"1ec187c9",
   819 => x"ddf64973",
   820 => x"c386c487",
   821 => x"731eecfe",
   822 => x"87f1f749",
   823 => x"4a6c86c4",
   824 => x"c404aa6d",
   825 => x"cf48ff87",
   826 => x"7ca2c187",
   827 => x"ffc74972",
   828 => x"ecfec399",
   829 => x"48699781",
   830 => x"4c264d26",
   831 => x"4f264b26",
   832 => x"711e731e",
   833 => x"c0029b4b",
   834 => x"cbc487e4",
   835 => x"4a735bdc",
   836 => x"c6c48ac2",
   837 => x"9249bfec",
   838 => x"bfc8cbc4",
   839 => x"c4807248",
   840 => x"7158e0cb",
   841 => x"c430c448",
   842 => x"c058fcc6",
   843 => x"cbc487ed",
   844 => x"cbc448d8",
   845 => x"c478bfcc",
   846 => x"c448dccb",
   847 => x"78bfd0cb",
   848 => x"bff4c6c4",
   849 => x"c487c902",
   850 => x"49bfecc6",
   851 => x"87c731c4",
   852 => x"bfd4cbc4",
   853 => x"c431c449",
   854 => x"2659fcc6",
   855 => x"0e4f264b",
   856 => x"0e5c5b5e",
   857 => x"4bc04a71",
   858 => x"c0029a72",
   859 => x"a2da87e1",
   860 => x"4b699f49",
   861 => x"bff4c6c4",
   862 => x"d487cf02",
   863 => x"699f49a2",
   864 => x"ffc04c49",
   865 => x"34d09cff",
   866 => x"4cc087c2",
   867 => x"73b34974",
   868 => x"87ecfd49",
   869 => x"4b264c26",
   870 => x"5e0e4f26",
   871 => x"0e5d5c5b",
   872 => x"a6c886f0",
   873 => x"ffffcf59",
   874 => x"c04cf8ff",
   875 => x"0266c47e",
   876 => x"fec387d8",
   877 => x"78c048e8",
   878 => x"48e0fec3",
   879 => x"bfdccbc4",
   880 => x"e4fec378",
   881 => x"d8cbc448",
   882 => x"c7c478bf",
   883 => x"50c048c9",
   884 => x"bff8c6c4",
   885 => x"e8fec349",
   886 => x"aa714abf",
   887 => x"87ccc403",
   888 => x"99cf4972",
   889 => x"87eac005",
   890 => x"48d8fec0",
   891 => x"bfe0fec3",
   892 => x"ecfec378",
   893 => x"e0fec31e",
   894 => x"fec349bf",
   895 => x"a1c148e0",
   896 => x"ddff7178",
   897 => x"86c487fe",
   898 => x"48d4fec0",
   899 => x"78ecfec3",
   900 => x"fec087cc",
   901 => x"c048bfd4",
   902 => x"fec080e0",
   903 => x"fec358d8",
   904 => x"c148bfe8",
   905 => x"ecfec380",
   906 => x"0f942758",
   907 => x"97bf0000",
   908 => x"029d4dbf",
   909 => x"c387e5c2",
   910 => x"c202ade5",
   911 => x"fec087de",
   912 => x"cb4bbfd4",
   913 => x"4c1149a3",
   914 => x"c105accf",
   915 => x"497587d2",
   916 => x"89c199df",
   917 => x"c6c491cd",
   918 => x"a3c181fc",
   919 => x"c351124a",
   920 => x"51124aa3",
   921 => x"124aa3c5",
   922 => x"4aa3c751",
   923 => x"a3c95112",
   924 => x"ce51124a",
   925 => x"51124aa3",
   926 => x"124aa3d0",
   927 => x"4aa3d251",
   928 => x"a3d45112",
   929 => x"d651124a",
   930 => x"51124aa3",
   931 => x"124aa3d8",
   932 => x"4aa3dc51",
   933 => x"a3de5112",
   934 => x"c151124a",
   935 => x"87fcc07e",
   936 => x"99c84974",
   937 => x"87edc005",
   938 => x"99d04974",
   939 => x"c087d305",
   940 => x"c00266e0",
   941 => x"497387cc",
   942 => x"0f66e0c0",
   943 => x"c0029870",
   944 => x"056e87d3",
   945 => x"c487c6c0",
   946 => x"c048fcc6",
   947 => x"d4fec050",
   948 => x"edc248bf",
   949 => x"c9c7c487",
   950 => x"7e50c048",
   951 => x"bff8c6c4",
   952 => x"e8fec349",
   953 => x"aa714abf",
   954 => x"87f4fb04",
   955 => x"ffffffcf",
   956 => x"cbc44cf8",
   957 => x"c005bfdc",
   958 => x"c6c487c8",
   959 => x"c102bff4",
   960 => x"fec387fe",
   961 => x"e849bfe4",
   962 => x"497087c6",
   963 => x"59e8fec3",
   964 => x"c348a6c4",
   965 => x"78bfe4fe",
   966 => x"bff4c6c4",
   967 => x"87dbc002",
   968 => x"744966c4",
   969 => x"02a97499",
   970 => x"c887c8c0",
   971 => x"78c048a6",
   972 => x"c887e7c0",
   973 => x"78c148a6",
   974 => x"c487dfc0",
   975 => x"ffcf4966",
   976 => x"02a999f8",
   977 => x"cc87c8c0",
   978 => x"78c048a6",
   979 => x"cc87c5c0",
   980 => x"78c148a6",
   981 => x"cc48a6c8",
   982 => x"66c87866",
   983 => x"87e0c005",
   984 => x"c24966c4",
   985 => x"ecc6c489",
   986 => x"c4914abf",
   987 => x"4abfc8cb",
   988 => x"48e0fec3",
   989 => x"c378a172",
   990 => x"c048e8fe",
   991 => x"87d0f978",
   992 => x"ffcf48c0",
   993 => x"4cf8ffff",
   994 => x"4d268ef0",
   995 => x"4b264c26",
   996 => x"00004f26",
   997 => x"00000000",
   998 => x"ffffffff",
   999 => x"00000fa4",
  1000 => x"00000fb0",
  1001 => x"33544146",
  1002 => x"20202032",
  1003 => x"00000000",
  1004 => x"31544146",
  1005 => x"20202036",
  1006 => x"d4ff1e00",
  1007 => x"78ffc348",
  1008 => x"4f264868",
  1009 => x"48d4ff1e",
  1010 => x"ff78ffc3",
  1011 => x"e1c048d0",
  1012 => x"48d4ff78",
  1013 => x"cbc478d4",
  1014 => x"d4ff48e0",
  1015 => x"4f2650bf",
  1016 => x"48d0ff1e",
  1017 => x"2678e0c0",
  1018 => x"ccff1e4f",
  1019 => x"99497087",
  1020 => x"c087c602",
  1021 => x"f105a9fb",
  1022 => x"26487187",
  1023 => x"5b5e0e4f",
  1024 => x"4b710e5c",
  1025 => x"f0fe4cc0",
  1026 => x"99497087",
  1027 => x"87f9c002",
  1028 => x"02a9ecc0",
  1029 => x"c087f2c0",
  1030 => x"c002a9fb",
  1031 => x"66cc87eb",
  1032 => x"c703acb7",
  1033 => x"0266d087",
  1034 => x"537187c2",
  1035 => x"c2029971",
  1036 => x"fe84c187",
  1037 => x"497087c3",
  1038 => x"87cd0299",
  1039 => x"02a9ecc0",
  1040 => x"fbc087c7",
  1041 => x"d5ff05a9",
  1042 => x"0266d087",
  1043 => x"97c087c3",
  1044 => x"a9ecc07b",
  1045 => x"7487c405",
  1046 => x"7487c54a",
  1047 => x"8a0ac04a",
  1048 => x"4c264872",
  1049 => x"4f264b26",
  1050 => x"87cdfd1e",
  1051 => x"c04a4970",
  1052 => x"c904aaf0",
  1053 => x"aaf9c087",
  1054 => x"c087c301",
  1055 => x"c1c18af0",
  1056 => x"87c904aa",
  1057 => x"01aadac1",
  1058 => x"f7c087c3",
  1059 => x"2648728a",
  1060 => x"5b5e0e4f",
  1061 => x"4a710e5c",
  1062 => x"724cd4ff",
  1063 => x"87ecc049",
  1064 => x"029b4b70",
  1065 => x"8bc187c2",
  1066 => x"c548d0ff",
  1067 => x"7cd5c178",
  1068 => x"31c64973",
  1069 => x"97dcf2c1",
  1070 => x"71484abf",
  1071 => x"ff7c70b0",
  1072 => x"78c448d0",
  1073 => x"4c264873",
  1074 => x"4f264b26",
  1075 => x"5c5b5e0e",
  1076 => x"86f80e5d",
  1077 => x"a6c44d71",
  1078 => x"fb78c048",
  1079 => x"4bc087e6",
  1080 => x"97ccc6c1",
  1081 => x"a9c049bf",
  1082 => x"fb87cf04",
  1083 => x"83c187fb",
  1084 => x"97ccc6c1",
  1085 => x"06ab49bf",
  1086 => x"c6c187f1",
  1087 => x"02bf97cc",
  1088 => x"f4fa87cf",
  1089 => x"99497087",
  1090 => x"c087c602",
  1091 => x"f105a9ec",
  1092 => x"754bc087",
  1093 => x"87e1fa7e",
  1094 => x"dcfa4c70",
  1095 => x"fa4d7087",
  1096 => x"4a7087d7",
  1097 => x"496e83c1",
  1098 => x"699781c8",
  1099 => x"c702ac49",
  1100 => x"acffc087",
  1101 => x"87e9c005",
  1102 => x"81c9496e",
  1103 => x"ad496997",
  1104 => x"c087c602",
  1105 => x"d805adff",
  1106 => x"ca496e87",
  1107 => x"49699781",
  1108 => x"87c602aa",
  1109 => x"05aaffc0",
  1110 => x"a6c487c7",
  1111 => x"d378c148",
  1112 => x"acecc087",
  1113 => x"c087c602",
  1114 => x"c705acfb",
  1115 => x"c44bc087",
  1116 => x"78c148a6",
  1117 => x"fe0266c4",
  1118 => x"e3f987db",
  1119 => x"f8487387",
  1120 => x"264d268e",
  1121 => x"264b264c",
  1122 => x"0000004f",
  1123 => x"5b5e0e00",
  1124 => x"f80e5d5c",
  1125 => x"ff7e7186",
  1126 => x"1e6e4bd4",
  1127 => x"49e8cbc4",
  1128 => x"87e3dfff",
  1129 => x"987086c4",
  1130 => x"87d0c402",
  1131 => x"c148a6c4",
  1132 => x"78bfe4f2",
  1133 => x"d8fb496e",
  1134 => x"48d0ff87",
  1135 => x"d6c178c5",
  1136 => x"6e4ac07b",
  1137 => x"11817249",
  1138 => x"cb82c17b",
  1139 => x"f204aab7",
  1140 => x"c34acc87",
  1141 => x"82c17bff",
  1142 => x"aab7e0c0",
  1143 => x"ff87f404",
  1144 => x"78c448d0",
  1145 => x"c57bffc3",
  1146 => x"7bd3c178",
  1147 => x"78c47bc1",
  1148 => x"66c47e73",
  1149 => x"a8b7c048",
  1150 => x"87eec206",
  1151 => x"bff0cbc4",
  1152 => x"4866c44c",
  1153 => x"a6c88874",
  1154 => x"029c7458",
  1155 => x"c387f7c1",
  1156 => x"c84decfe",
  1157 => x"c08c4bc0",
  1158 => x"c603acb7",
  1159 => x"a4c0c887",
  1160 => x"c44cc04b",
  1161 => x"bf97e0cb",
  1162 => x"0299d049",
  1163 => x"1ec087d1",
  1164 => x"49e8cbc4",
  1165 => x"c487d6e2",
  1166 => x"4a497086",
  1167 => x"c387ebc0",
  1168 => x"c41eecfe",
  1169 => x"e249e8cb",
  1170 => x"86c487c3",
  1171 => x"ff4a4970",
  1172 => x"c5c848d0",
  1173 => x"c1486e78",
  1174 => x"481578d4",
  1175 => x"c178086e",
  1176 => x"f5ff058b",
  1177 => x"48d0ff87",
  1178 => x"9a7278c4",
  1179 => x"c087c505",
  1180 => x"87cac148",
  1181 => x"cbc41ec1",
  1182 => x"dfff49e8",
  1183 => x"86c487f0",
  1184 => x"fe059c74",
  1185 => x"66c487c9",
  1186 => x"a8b7c048",
  1187 => x"c487d106",
  1188 => x"c048e8cb",
  1189 => x"c080d078",
  1190 => x"c480f478",
  1191 => x"78bff4cb",
  1192 => x"c04866c4",
  1193 => x"fd01a8b7",
  1194 => x"4b6e87d2",
  1195 => x"c548d0ff",
  1196 => x"7bd3c178",
  1197 => x"78c47bc0",
  1198 => x"87c248c1",
  1199 => x"8ef848c0",
  1200 => x"4c264d26",
  1201 => x"4f264b26",
  1202 => x"5c5b5e0e",
  1203 => x"86fc0e5d",
  1204 => x"4bc04d71",
  1205 => x"c004ad4c",
  1206 => x"c3c187e8",
  1207 => x"9c741ecc",
  1208 => x"c087c402",
  1209 => x"c187c24a",
  1210 => x"ea49724a",
  1211 => x"86c487ec",
  1212 => x"83c17e70",
  1213 => x"87c2056e",
  1214 => x"84c14b75",
  1215 => x"ff06ab75",
  1216 => x"486e87d8",
  1217 => x"4d268efc",
  1218 => x"4b264c26",
  1219 => x"711e4f26",
  1220 => x"ffc3494a",
  1221 => x"48d4ff99",
  1222 => x"49727871",
  1223 => x"c329b7c8",
  1224 => x"787199ff",
  1225 => x"b7d04972",
  1226 => x"99ffc329",
  1227 => x"49727871",
  1228 => x"c329b7d8",
  1229 => x"787199ff",
  1230 => x"5e0e4f26",
  1231 => x"0e5d5c5b",
  1232 => x"4a7186fc",
  1233 => x"49724cc0",
  1234 => x"87ffecc1",
  1235 => x"da059870",
  1236 => x"734bc187",
  1237 => x"d2eec149",
  1238 => x"05987087",
  1239 => x"4cc187c2",
  1240 => x"d1c483c1",
  1241 => x"abb7bfc4",
  1242 => x"ff87e806",
  1243 => x"e1c848d0",
  1244 => x"48d4ff78",
  1245 => x"9c7478dd",
  1246 => x"c487c702",
  1247 => x"4dbfecd1",
  1248 => x"4dc087c2",
  1249 => x"c5fe4975",
  1250 => x"029c7487",
  1251 => x"d1c487c7",
  1252 => x"c27ebfec",
  1253 => x"6e7ec087",
  1254 => x"87f2fd49",
  1255 => x"edfd49c0",
  1256 => x"fd49c087",
  1257 => x"d0ff87e8",
  1258 => x"78e0c048",
  1259 => x"49dc1ec1",
  1260 => x"87dafbc0",
  1261 => x"8ef84874",
  1262 => x"4c264d26",
  1263 => x"4f264b26",
  1264 => x"c44a711e",
  1265 => x"87c90266",
  1266 => x"89c3c149",
  1267 => x"cc87c902",
  1268 => x"f6497287",
  1269 => x"87c587f7",
  1270 => x"ddfd4972",
  1271 => x"0e4f2687",
  1272 => x"5d5c5b5e",
  1273 => x"7186fc0e",
  1274 => x"91de494c",
  1275 => x"4dd0ccc4",
  1276 => x"6d978571",
  1277 => x"87dcc102",
  1278 => x"bffccbc4",
  1279 => x"7282744a",
  1280 => x"87c4fb49",
  1281 => x"026e7e70",
  1282 => x"c487f2c0",
  1283 => x"6e4bc4cc",
  1284 => x"fe49cb4a",
  1285 => x"7487e2f2",
  1286 => x"c193cc4b",
  1287 => x"c483f8f2",
  1288 => x"e0d1c183",
  1289 => x"c149747b",
  1290 => x"7587d1cd",
  1291 => x"e0f2c17b",
  1292 => x"1e49bf97",
  1293 => x"49c4ccc4",
  1294 => x"c487c5fe",
  1295 => x"c1497486",
  1296 => x"c087f9cc",
  1297 => x"d4cec149",
  1298 => x"e4cbc487",
  1299 => x"c178c048",
  1300 => x"87efdd49",
  1301 => x"4d268efc",
  1302 => x"4b264c26",
  1303 => x"00004f26",
  1304 => x"64616f4c",
  1305 => x"2e676e69",
  1306 => x"0e002e2e",
  1307 => x"0e5c5b5e",
  1308 => x"c44a4b71",
  1309 => x"82bffccb",
  1310 => x"cbf94972",
  1311 => x"9c4c7087",
  1312 => x"4987c402",
  1313 => x"c487d8e3",
  1314 => x"c048fccb",
  1315 => x"dc49c178",
  1316 => x"4c2687f1",
  1317 => x"4f264b26",
  1318 => x"5c5b5e0e",
  1319 => x"86f40e5d",
  1320 => x"4decfec3",
  1321 => x"a6c44cc0",
  1322 => x"c478c048",
  1323 => x"49bffccb",
  1324 => x"a9c07e75",
  1325 => x"87fbc006",
  1326 => x"fec37e75",
  1327 => x"029848ec",
  1328 => x"c187f0c0",
  1329 => x"c81eccc3",
  1330 => x"87c40266",
  1331 => x"87c24dc0",
  1332 => x"49754dc1",
  1333 => x"c487c3e3",
  1334 => x"c17e7086",
  1335 => x"4866c484",
  1336 => x"a6c880c1",
  1337 => x"fccbc458",
  1338 => x"03ac49bf",
  1339 => x"056e87c5",
  1340 => x"6e87d0ff",
  1341 => x"754cc04d",
  1342 => x"e0c3029d",
  1343 => x"ccc3c187",
  1344 => x"0266c81e",
  1345 => x"a6cc87c7",
  1346 => x"c578c048",
  1347 => x"48a6cc87",
  1348 => x"66cc78c1",
  1349 => x"87c2e249",
  1350 => x"7e7086c4",
  1351 => x"e9c2026e",
  1352 => x"cb496e87",
  1353 => x"49699781",
  1354 => x"c10299d0",
  1355 => x"d1c187d6",
  1356 => x"49744aeb",
  1357 => x"f2c191cc",
  1358 => x"797281f8",
  1359 => x"ffc381c8",
  1360 => x"de497451",
  1361 => x"d0ccc491",
  1362 => x"c285714d",
  1363 => x"c17d97c1",
  1364 => x"e0c049a5",
  1365 => x"fcc6c451",
  1366 => x"d202bf97",
  1367 => x"c284c187",
  1368 => x"c6c44ba5",
  1369 => x"49db4afc",
  1370 => x"87cdedfe",
  1371 => x"cd87dbc1",
  1372 => x"51c049a5",
  1373 => x"a5c284c1",
  1374 => x"cb4a6e4b",
  1375 => x"f8ecfe49",
  1376 => x"87c6c187",
  1377 => x"4adfcfc1",
  1378 => x"91cc4974",
  1379 => x"81f8f2c1",
  1380 => x"c6c47972",
  1381 => x"02bf97fc",
  1382 => x"497487d8",
  1383 => x"84c191de",
  1384 => x"4bd0ccc4",
  1385 => x"c6c48371",
  1386 => x"49dd4afc",
  1387 => x"87c9ecfe",
  1388 => x"4b7487d8",
  1389 => x"ccc493de",
  1390 => x"a3cb83d0",
  1391 => x"c151c049",
  1392 => x"4a6e7384",
  1393 => x"ebfe49cb",
  1394 => x"66c487ef",
  1395 => x"c880c148",
  1396 => x"acc758a6",
  1397 => x"87c5c003",
  1398 => x"e0fc056e",
  1399 => x"f4487487",
  1400 => x"264d268e",
  1401 => x"264b264c",
  1402 => x"1e731e4f",
  1403 => x"cc494b71",
  1404 => x"f8f2c191",
  1405 => x"4aa1c881",
  1406 => x"48dcf2c1",
  1407 => x"a1c95012",
  1408 => x"ccc6c14a",
  1409 => x"ca501248",
  1410 => x"e0f2c181",
  1411 => x"c1501148",
  1412 => x"bf97e0f2",
  1413 => x"49c01e49",
  1414 => x"c487e5f6",
  1415 => x"de48e4cb",
  1416 => x"d649c178",
  1417 => x"8efc87dd",
  1418 => x"4f264b26",
  1419 => x"494a711e",
  1420 => x"f2c191cc",
  1421 => x"81c881f8",
  1422 => x"cbc44811",
  1423 => x"cbc458e8",
  1424 => x"78c048fc",
  1425 => x"fad549c1",
  1426 => x"1e4f2687",
  1427 => x"c6c149c0",
  1428 => x"4f2687cb",
  1429 => x"0299711e",
  1430 => x"f4c187d2",
  1431 => x"50c048d4",
  1432 => x"d8c180f7",
  1433 => x"f2c140ec",
  1434 => x"87ce78f0",
  1435 => x"48d0f4c1",
  1436 => x"78e8f2c1",
  1437 => x"d9c180fc",
  1438 => x"4f2678cb",
  1439 => x"5c5b5e0e",
  1440 => x"4a4c710e",
  1441 => x"f2c192cc",
  1442 => x"a2c882f8",
  1443 => x"4ba2c949",
  1444 => x"1e4b6b97",
  1445 => x"1e496997",
  1446 => x"491282ca",
  1447 => x"87caf1c0",
  1448 => x"ded449c0",
  1449 => x"c1497487",
  1450 => x"f887d1c3",
  1451 => x"264c268e",
  1452 => x"1e4f264b",
  1453 => x"4b711e73",
  1454 => x"87c0ff49",
  1455 => x"fbfe4973",
  1456 => x"264b2687",
  1457 => x"1e731e4f",
  1458 => x"a3c64b71",
  1459 => x"87db024a",
  1460 => x"d6028ac1",
  1461 => x"c1028a87",
  1462 => x"028a87da",
  1463 => x"8a87fcc0",
  1464 => x"87e1c002",
  1465 => x"87cb028a",
  1466 => x"c787dbc1",
  1467 => x"87fcfc49",
  1468 => x"c487dec1",
  1469 => x"02bffccb",
  1470 => x"4887cbc1",
  1471 => x"ccc488c1",
  1472 => x"c1c158c0",
  1473 => x"c0ccc487",
  1474 => x"f9c002bf",
  1475 => x"fccbc487",
  1476 => x"80c148bf",
  1477 => x"58c0ccc4",
  1478 => x"c487ebc0",
  1479 => x"49bffccb",
  1480 => x"ccc489c6",
  1481 => x"b7c059c0",
  1482 => x"87da03a9",
  1483 => x"48fccbc4",
  1484 => x"87d278c0",
  1485 => x"bfc0ccc4",
  1486 => x"c487cb02",
  1487 => x"48bffccb",
  1488 => x"ccc480c6",
  1489 => x"49c058c0",
  1490 => x"7387f8d1",
  1491 => x"ebc0c149",
  1492 => x"264b2687",
  1493 => x"5b5e0e4f",
  1494 => x"ff0e5d5c",
  1495 => x"a6dc86d0",
  1496 => x"48a6c859",
  1497 => x"80c478c0",
  1498 => x"7866c4c1",
  1499 => x"78c180c4",
  1500 => x"78c180c4",
  1501 => x"48c0ccc4",
  1502 => x"cbc478c1",
  1503 => x"de48bfe4",
  1504 => x"87cb05a8",
  1505 => x"7087d1f4",
  1506 => x"59a6cc49",
  1507 => x"e087edcf",
  1508 => x"d4e187f2",
  1509 => x"87e1e087",
  1510 => x"fbc04c70",
  1511 => x"f1c102ac",
  1512 => x"0566d887",
  1513 => x"c187e2c1",
  1514 => x"c44a66c0",
  1515 => x"c17e6a82",
  1516 => x"6e48f4ee",
  1517 => x"20412049",
  1518 => x"c1511041",
  1519 => x"c14866c0",
  1520 => x"6a78e9d7",
  1521 => x"7481c749",
  1522 => x"66c0c151",
  1523 => x"c181c849",
  1524 => x"66c0c151",
  1525 => x"c081c949",
  1526 => x"66c0c151",
  1527 => x"c081ca49",
  1528 => x"d81ec151",
  1529 => x"c8496a1e",
  1530 => x"87d1e081",
  1531 => x"c4c186c8",
  1532 => x"a8c04866",
  1533 => x"c887c701",
  1534 => x"78c148a6",
  1535 => x"c4c187cf",
  1536 => x"88c14866",
  1537 => x"c458a6d0",
  1538 => x"dcdfff87",
  1539 => x"48a6d087",
  1540 => x"9c7478c2",
  1541 => x"87e0cd02",
  1542 => x"c14866c8",
  1543 => x"03a866c8",
  1544 => x"dc87d5cd",
  1545 => x"78c048a6",
  1546 => x"ccdeff7e",
  1547 => x"c14c7087",
  1548 => x"c205acd0",
  1549 => x"a6c487da",
  1550 => x"e0786e48",
  1551 => x"497087ea",
  1552 => x"f4ddff7e",
  1553 => x"c04c7087",
  1554 => x"c105acec",
  1555 => x"66c887ed",
  1556 => x"c191cc49",
  1557 => x"c48166c0",
  1558 => x"4d6a4aa1",
  1559 => x"6e4aa1c8",
  1560 => x"ecd8c152",
  1561 => x"d0ddff79",
  1562 => x"9c4c7087",
  1563 => x"c087d902",
  1564 => x"d302acfb",
  1565 => x"ff557487",
  1566 => x"7087fedc",
  1567 => x"c7029c4c",
  1568 => x"acfbc087",
  1569 => x"87edff05",
  1570 => x"c255e0c0",
  1571 => x"97c055c1",
  1572 => x"4966d87d",
  1573 => x"05a966c4",
  1574 => x"66c887db",
  1575 => x"a866cc48",
  1576 => x"c887ca04",
  1577 => x"80c14866",
  1578 => x"c858a6cc",
  1579 => x"4866cc87",
  1580 => x"a6d088c1",
  1581 => x"c0dcff58",
  1582 => x"c14c7087",
  1583 => x"c805acd0",
  1584 => x"4866d487",
  1585 => x"a6d880c1",
  1586 => x"acd0c158",
  1587 => x"87e6fd02",
  1588 => x"48a6e0c0",
  1589 => x"6e7866d8",
  1590 => x"66e0c048",
  1591 => x"e9c905a8",
  1592 => x"a6e4c087",
  1593 => x"e078c048",
  1594 => x"7478c080",
  1595 => x"88fbc048",
  1596 => x"58a6ecc0",
  1597 => x"c8029870",
  1598 => x"cb4887ea",
  1599 => x"a6ecc088",
  1600 => x"02987058",
  1601 => x"4887d3c1",
  1602 => x"ecc088c9",
  1603 => x"987058a6",
  1604 => x"87edc302",
  1605 => x"c088c448",
  1606 => x"7058a6ec",
  1607 => x"87d00298",
  1608 => x"c088c148",
  1609 => x"7058a6ec",
  1610 => x"d4c30298",
  1611 => x"87eec787",
  1612 => x"c048a6dc",
  1613 => x"d9ff78f0",
  1614 => x"4c7087ff",
  1615 => x"02acecc0",
  1616 => x"c087c4c0",
  1617 => x"c05ca6e0",
  1618 => x"cd02acec",
  1619 => x"e8d9ff87",
  1620 => x"c04c7087",
  1621 => x"ff05acec",
  1622 => x"ecc087f3",
  1623 => x"c4c002ac",
  1624 => x"d4d9ff87",
  1625 => x"ca1ec087",
  1626 => x"4966d01e",
  1627 => x"c8c191cc",
  1628 => x"80714866",
  1629 => x"c858a6cc",
  1630 => x"80c44866",
  1631 => x"cc58a6d0",
  1632 => x"ff49bf66",
  1633 => x"c187f6d9",
  1634 => x"d41ede1e",
  1635 => x"ff49bf66",
  1636 => x"d087ead9",
  1637 => x"c0497086",
  1638 => x"ecc08909",
  1639 => x"e8c059a6",
  1640 => x"a8c04866",
  1641 => x"87eec006",
  1642 => x"4866e8c0",
  1643 => x"c003a8dd",
  1644 => x"66c487e4",
  1645 => x"e8c049bf",
  1646 => x"e0c08166",
  1647 => x"66e8c051",
  1648 => x"c481c149",
  1649 => x"c281bf66",
  1650 => x"e8c051c1",
  1651 => x"81c24966",
  1652 => x"81bf66c4",
  1653 => x"486e51c0",
  1654 => x"78e9d7c1",
  1655 => x"81c8496e",
  1656 => x"6e5166d0",
  1657 => x"d481c949",
  1658 => x"496e5166",
  1659 => x"66dc81ca",
  1660 => x"4866d051",
  1661 => x"a6d480c1",
  1662 => x"80f44858",
  1663 => x"e3c478c1",
  1664 => x"e3d9ff87",
  1665 => x"c0497087",
  1666 => x"ff59a6ec",
  1667 => x"7087d9d9",
  1668 => x"a6e0c049",
  1669 => x"4866dc59",
  1670 => x"05a8ecc0",
  1671 => x"dc87cac0",
  1672 => x"e8c048a6",
  1673 => x"c4c07866",
  1674 => x"ccd6ff87",
  1675 => x"4966c887",
  1676 => x"c0c191cc",
  1677 => x"80714866",
  1678 => x"c458a6c8",
  1679 => x"82c84a66",
  1680 => x"ca4966c4",
  1681 => x"66e8c081",
  1682 => x"4966dc51",
  1683 => x"e8c081c1",
  1684 => x"48c18966",
  1685 => x"49703071",
  1686 => x"977189c1",
  1687 => x"d4d0c47a",
  1688 => x"e8c049bf",
  1689 => x"6a972966",
  1690 => x"9871484a",
  1691 => x"58a6f0c0",
  1692 => x"c44966c4",
  1693 => x"c04d6981",
  1694 => x"6e4866e0",
  1695 => x"c5c002a8",
  1696 => x"c07ec087",
  1697 => x"7ec187c2",
  1698 => x"e0c01e6e",
  1699 => x"ff49751e",
  1700 => x"c887ead5",
  1701 => x"c04c7086",
  1702 => x"c106acb7",
  1703 => x"857487d0",
  1704 => x"7449e0c0",
  1705 => x"c14b7589",
  1706 => x"714ac0ef",
  1707 => x"87c9d8fe",
  1708 => x"7e7585c2",
  1709 => x"4866e4c0",
  1710 => x"e8c080c1",
  1711 => x"ecc058a6",
  1712 => x"81c14966",
  1713 => x"c002a970",
  1714 => x"4dc087c5",
  1715 => x"c187c2c0",
  1716 => x"c21e754d",
  1717 => x"e0c049a4",
  1718 => x"70887148",
  1719 => x"66c81e49",
  1720 => x"d8d4ff49",
  1721 => x"c086c887",
  1722 => x"ff01a8b7",
  1723 => x"e4c087c6",
  1724 => x"d3c00266",
  1725 => x"4966c487",
  1726 => x"e4c081c9",
  1727 => x"66c45166",
  1728 => x"fcd9c148",
  1729 => x"87cec078",
  1730 => x"c94966c4",
  1731 => x"c451c281",
  1732 => x"dac14866",
  1733 => x"a6c478f3",
  1734 => x"c078c148",
  1735 => x"d3ff87c6",
  1736 => x"4c7087c7",
  1737 => x"c00266c4",
  1738 => x"66c887f5",
  1739 => x"a866cc48",
  1740 => x"87cbc004",
  1741 => x"c14866c8",
  1742 => x"58a6cc80",
  1743 => x"cc87e0c0",
  1744 => x"88c14866",
  1745 => x"c058a6d0",
  1746 => x"c6c187d5",
  1747 => x"c8c005ac",
  1748 => x"4866d087",
  1749 => x"a6d480c1",
  1750 => x"ccd2ff58",
  1751 => x"d44c7087",
  1752 => x"80c14866",
  1753 => x"7458a6d8",
  1754 => x"cbc0029c",
  1755 => x"4866c887",
  1756 => x"a866c8c1",
  1757 => x"87ebf204",
  1758 => x"87e4d1ff",
  1759 => x"c74866c8",
  1760 => x"e1c003a8",
  1761 => x"4c66c887",
  1762 => x"48c0ccc4",
  1763 => x"497478c0",
  1764 => x"c0c191cc",
  1765 => x"a1c48166",
  1766 => x"c04a6a4a",
  1767 => x"84c17952",
  1768 => x"ff04acc7",
  1769 => x"d0ff87e2",
  1770 => x"264d268e",
  1771 => x"264b264c",
  1772 => x"0000004f",
  1773 => x"64616f4c",
  1774 => x"202e2a20",
  1775 => x"00000000",
  1776 => x"1e00203a",
  1777 => x"4b711e73",
  1778 => x"87c6029b",
  1779 => x"48fccbc4",
  1780 => x"1ec778c0",
  1781 => x"bffccbc4",
  1782 => x"f2c11e49",
  1783 => x"cbc41ef8",
  1784 => x"ed49bfe4",
  1785 => x"86cc87ef",
  1786 => x"bfe4cbc4",
  1787 => x"87e4e949",
  1788 => x"c8029b73",
  1789 => x"f8f2c187",
  1790 => x"cdefc049",
  1791 => x"264b2687",
  1792 => x"eccc1e4f",
  1793 => x"fe49c187",
  1794 => x"e2fe87f9",
  1795 => x"987087d7",
  1796 => x"fe87cd02",
  1797 => x"7087fee9",
  1798 => x"87c40298",
  1799 => x"87c24ac1",
  1800 => x"9a724ac0",
  1801 => x"c087ce05",
  1802 => x"d8f1c11e",
  1803 => x"d1fcc049",
  1804 => x"fe86c487",
  1805 => x"e5cbc287",
  1806 => x"c11ec087",
  1807 => x"c049e4f1",
  1808 => x"c087fffb",
  1809 => x"ffcbc21e",
  1810 => x"c0497087",
  1811 => x"c387f3fb",
  1812 => x"8ef887ea",
  1813 => x"00004f26",
  1814 => x"66204453",
  1815 => x"656c6961",
  1816 => x"00002e64",
  1817 => x"746f6f42",
  1818 => x"2e676e69",
  1819 => x"1e002e2e",
  1820 => x"e7d049c0",
  1821 => x"edc6c287",
  1822 => x"f6f1c087",
  1823 => x"e5c6c287",
  1824 => x"2687ed87",
  1825 => x"cbc41e4f",
  1826 => x"78c048fc",
  1827 => x"48e4cbc4",
  1828 => x"ecfd78c0",
  1829 => x"87d7ff87",
  1830 => x"4f2648c0",
  1831 => x"00000000",
  1832 => x"00000000",
  1833 => x"00000001",
  1834 => x"78452080",
  1835 => x"00007469",
  1836 => x"61422080",
  1837 => x"00006b63",
  1838 => x"0000162c",
  1839 => x"00004310",
  1840 => x"00000000",
  1841 => x"0000162c",
  1842 => x"0000432e",
  1843 => x"00000000",
  1844 => x"0000162c",
  1845 => x"0000434c",
  1846 => x"00000000",
  1847 => x"0000162c",
  1848 => x"0000436a",
  1849 => x"00000000",
  1850 => x"0000162c",
  1851 => x"00004388",
  1852 => x"00000000",
  1853 => x"0000162c",
  1854 => x"000043a6",
  1855 => x"00000000",
  1856 => x"0000162c",
  1857 => x"000043c4",
  1858 => x"00000000",
  1859 => x"0000162c",
  1860 => x"00000000",
  1861 => x"00000000",
  1862 => x"000016c5",
  1863 => x"00000000",
  1864 => x"00000000",
  1865 => x"48f0fe1e",
  1866 => x"09cd78c0",
  1867 => x"4f260979",
  1868 => x"fe86fc1e",
  1869 => x"487ebff0",
  1870 => x"4f268efc",
  1871 => x"48f0fe1e",
  1872 => x"4f2678c1",
  1873 => x"48f0fe1e",
  1874 => x"4f2678c0",
  1875 => x"c04a711e",
  1876 => x"a2c17a97",
  1877 => x"ca51c049",
  1878 => x"51c049a2",
  1879 => x"c049a2cb",
  1880 => x"0e4f2651",
  1881 => x"0e5c5b5e",
  1882 => x"4c7186f0",
  1883 => x"9749a4ca",
  1884 => x"a4cb7e69",
  1885 => x"486b974b",
  1886 => x"c158a6c8",
  1887 => x"58a6cc80",
  1888 => x"a6d098c7",
  1889 => x"cc486e58",
  1890 => x"db05a866",
  1891 => x"7e699787",
  1892 => x"c8486b97",
  1893 => x"80c158a6",
  1894 => x"c758a6cc",
  1895 => x"58a6d098",
  1896 => x"66cc486e",
  1897 => x"87e502a8",
  1898 => x"cc87d9fe",
  1899 => x"6b974aa4",
  1900 => x"49a17249",
  1901 => x"975166dc",
  1902 => x"486e7e6b",
  1903 => x"a6c880c1",
  1904 => x"cc98c758",
  1905 => x"977058a6",
  1906 => x"87d1c27b",
  1907 => x"f087edfd",
  1908 => x"264c268e",
  1909 => x"0e4f264b",
  1910 => x"5d5c5b5e",
  1911 => x"7186f40e",
  1912 => x"7e6d974d",
  1913 => x"974ca5c1",
  1914 => x"a6c8486c",
  1915 => x"c4486e58",
  1916 => x"c505a866",
  1917 => x"c048ff87",
  1918 => x"c7fd87e6",
  1919 => x"49a5c287",
  1920 => x"714b6c97",
  1921 => x"6b974ba3",
  1922 => x"7e6c974b",
  1923 => x"80c1486e",
  1924 => x"c758a6c8",
  1925 => x"58a6cc98",
  1926 => x"fc7c9770",
  1927 => x"487387de",
  1928 => x"4d268ef4",
  1929 => x"4b264c26",
  1930 => x"5e0e4f26",
  1931 => x"f40e5c5b",
  1932 => x"d84c7186",
  1933 => x"ffc34a66",
  1934 => x"4ba4c29a",
  1935 => x"73496c97",
  1936 => x"517249a1",
  1937 => x"6e7e6c97",
  1938 => x"c880c148",
  1939 => x"98c758a6",
  1940 => x"7058a6cc",
  1941 => x"268ef454",
  1942 => x"264b264c",
  1943 => x"1e731e4f",
  1944 => x"dffb86f4",
  1945 => x"4bbfe087",
  1946 => x"c0e0c049",
  1947 => x"87cb0299",
  1948 => x"cfc41e73",
  1949 => x"f1fe49e4",
  1950 => x"7386c487",
  1951 => x"99c0d049",
  1952 => x"87c0c102",
  1953 => x"97eecfc4",
  1954 => x"cfc47ebf",
  1955 => x"48bf97ef",
  1956 => x"6e58a6c8",
  1957 => x"a866c448",
  1958 => x"87e8c002",
  1959 => x"97eecfc4",
  1960 => x"cfc449bf",
  1961 => x"481181f0",
  1962 => x"c47808e0",
  1963 => x"bf97eecf",
  1964 => x"c1486e7e",
  1965 => x"58a6c880",
  1966 => x"a6cc98c7",
  1967 => x"eecfc458",
  1968 => x"5066c848",
  1969 => x"494bbfe4",
  1970 => x"99c0e0c0",
  1971 => x"7387cb02",
  1972 => x"f8cfc41e",
  1973 => x"87d2fd49",
  1974 => x"497386c4",
  1975 => x"0299c0d0",
  1976 => x"c487c0c1",
  1977 => x"bf97c2d0",
  1978 => x"c3d0c47e",
  1979 => x"c848bf97",
  1980 => x"486e58a6",
  1981 => x"02a866c4",
  1982 => x"c487e8c0",
  1983 => x"bf97c2d0",
  1984 => x"c4d0c449",
  1985 => x"e4481181",
  1986 => x"d0c47808",
  1987 => x"7ebf97c2",
  1988 => x"80c1486e",
  1989 => x"c758a6c8",
  1990 => x"58a6cc98",
  1991 => x"48c2d0c4",
  1992 => x"f85066c8",
  1993 => x"7e7087ca",
  1994 => x"f487d1f8",
  1995 => x"264b268e",
  1996 => x"cfc41e4f",
  1997 => x"d3f849e4",
  1998 => x"f8cfc487",
  1999 => x"87ccf849",
  2000 => x"49ddf9c1",
  2001 => x"c287ddf7",
  2002 => x"4f2687fb",
  2003 => x"c41e731e",
  2004 => x"fa49e4cf",
  2005 => x"4a7087c1",
  2006 => x"04aab7c0",
  2007 => x"c387ccc2",
  2008 => x"c905aaf0",
  2009 => x"f4ffc187",
  2010 => x"c178c148",
  2011 => x"e0c387ed",
  2012 => x"87c905aa",
  2013 => x"48f8ffc1",
  2014 => x"dec178c1",
  2015 => x"f8ffc187",
  2016 => x"87c602bf",
  2017 => x"4ba2c0c2",
  2018 => x"4b7287c2",
  2019 => x"bff4ffc1",
  2020 => x"87e0c002",
  2021 => x"b7c44973",
  2022 => x"c1c29129",
  2023 => x"4a7381dc",
  2024 => x"92c29acf",
  2025 => x"307248c1",
  2026 => x"baff4a70",
  2027 => x"98694872",
  2028 => x"87db7970",
  2029 => x"b7c44973",
  2030 => x"c1c29129",
  2031 => x"4a7381dc",
  2032 => x"92c29acf",
  2033 => x"307248c3",
  2034 => x"69484a70",
  2035 => x"c17970b0",
  2036 => x"c048f8ff",
  2037 => x"f4ffc178",
  2038 => x"c478c048",
  2039 => x"f749e4cf",
  2040 => x"4a7087f5",
  2041 => x"03aab7c0",
  2042 => x"c087f4fd",
  2043 => x"264b2648",
  2044 => x"0000004f",
  2045 => x"00000000",
  2046 => x"00000000",
  2047 => x"494a711e",
  2048 => x"2687c9fd",
  2049 => x"4ac01e4f",
  2050 => x"91c44972",
  2051 => x"81dcc1c2",
  2052 => x"82c179c0",
  2053 => x"04aab7d0",
  2054 => x"4f2687ee",
  2055 => x"5c5b5e0e",
  2056 => x"4d710e5d",
  2057 => x"7587ddf4",
  2058 => x"2ab7c44a",
  2059 => x"dcc1c292",
  2060 => x"cf4c7582",
  2061 => x"6a94c29c",
  2062 => x"2b744b49",
  2063 => x"48c29bc3",
  2064 => x"4c703074",
  2065 => x"4874bcff",
  2066 => x"7a709871",
  2067 => x"7387edf3",
  2068 => x"264d2648",
  2069 => x"264b264c",
  2070 => x"0000004f",
  2071 => x"00000000",
  2072 => x"00000000",
  2073 => x"00000000",
  2074 => x"00000000",
  2075 => x"00000000",
  2076 => x"00000000",
  2077 => x"00000000",
  2078 => x"00000000",
  2079 => x"00000000",
  2080 => x"00000000",
  2081 => x"00000000",
  2082 => x"00000000",
  2083 => x"00000000",
  2084 => x"00000000",
  2085 => x"00000000",
  2086 => x"00000000",
  2087 => x"5c5b5e0e",
  2088 => x"4a710e5d",
  2089 => x"724dd4ff",
  2090 => x"87c6029a",
  2091 => x"48d8c9c2",
  2092 => x"c9c278c0",
  2093 => x"c005bfd8",
  2094 => x"cfc487f9",
  2095 => x"d6f449f8",
  2096 => x"a8b7c087",
  2097 => x"c487cd04",
  2098 => x"f449f8cf",
  2099 => x"b7c087c9",
  2100 => x"87f303a8",
  2101 => x"bfd8c9c2",
  2102 => x"d8c9c249",
  2103 => x"78a1c148",
  2104 => x"81e8c9c2",
  2105 => x"c9c24811",
  2106 => x"c9c258e0",
  2107 => x"78c048e0",
  2108 => x"c287d8c5",
  2109 => x"02bfe0c9",
  2110 => x"c487f2c1",
  2111 => x"f349f8cf",
  2112 => x"b7c087d5",
  2113 => x"87cd04a8",
  2114 => x"bfe0c9c2",
  2115 => x"c288c148",
  2116 => x"db58e4c9",
  2117 => x"ccd0c487",
  2118 => x"f6c149bf",
  2119 => x"987087fe",
  2120 => x"c487cd02",
  2121 => x"f049f8cf",
  2122 => x"c9c287e2",
  2123 => x"78c048d8",
  2124 => x"bfdcc9c2",
  2125 => x"87d3c405",
  2126 => x"bfe0c9c2",
  2127 => x"87cbc405",
  2128 => x"bfd8c9c2",
  2129 => x"d8c9c249",
  2130 => x"78a1c148",
  2131 => x"81e8c9c2",
  2132 => x"c2494c11",
  2133 => x"c00299c0",
  2134 => x"487487cc",
  2135 => x"c298ffc1",
  2136 => x"c358e4c9",
  2137 => x"c9c287e5",
  2138 => x"dec35ce0",
  2139 => x"dcc9c287",
  2140 => x"ffc002bf",
  2141 => x"d8c9c287",
  2142 => x"c9c249bf",
  2143 => x"a1c148d8",
  2144 => x"e8c9c278",
  2145 => x"49699781",
  2146 => x"f8cfc41e",
  2147 => x"87d3ef49",
  2148 => x"c9c286c4",
  2149 => x"c148bfdc",
  2150 => x"e0c9c288",
  2151 => x"e0c9c258",
  2152 => x"c078c148",
  2153 => x"c149ecf6",
  2154 => x"7087e5f4",
  2155 => x"d0d0c449",
  2156 => x"87d7c259",
  2157 => x"49f8cfc4",
  2158 => x"7087dcf0",
  2159 => x"abb7c04b",
  2160 => x"87c7c204",
  2161 => x"bfd4c9c2",
  2162 => x"87e0c002",
  2163 => x"bfccd0c4",
  2164 => x"c7f4c149",
  2165 => x"02987087",
  2166 => x"c787d1c0",
  2167 => x"e4c9c248",
  2168 => x"c9c288bf",
  2169 => x"c9c258e8",
  2170 => x"78c048d4",
  2171 => x"bfd4c9c2",
  2172 => x"49a2c14a",
  2173 => x"59d8c9c2",
  2174 => x"82d0d0c4",
  2175 => x"c9c25273",
  2176 => x"a9b7bfe4",
  2177 => x"87e6c004",
  2178 => x"97d0d0c4",
  2179 => x"c41e49bf",
  2180 => x"87e4c149",
  2181 => x"d0c486c4",
  2182 => x"7dbf97d1",
  2183 => x"97d2d0c4",
  2184 => x"d0ff7dbf",
  2185 => x"78e0c048",
  2186 => x"48d4c9c2",
  2187 => x"f4c778c0",
  2188 => x"dbf2c149",
  2189 => x"c4497087",
  2190 => x"c459d0d0",
  2191 => x"ee49f8cf",
  2192 => x"4b7087d5",
  2193 => x"03abb7c0",
  2194 => x"2687f9fd",
  2195 => x"264c264d",
  2196 => x"004f264b",
  2197 => x"00000000",
  2198 => x"00000000",
  2199 => x"00000000",
  2200 => x"00000000",
  2201 => x"00000004",
  2202 => x"0882ff01",
  2203 => x"64f3c8f3",
  2204 => x"01f250f3",
  2205 => x"00f40181",
  2206 => x"48d0ff1e",
  2207 => x"7178e1c8",
  2208 => x"08d4ff48",
  2209 => x"4866c478",
  2210 => x"7808d4ff",
  2211 => x"711e4f26",
  2212 => x"4966c44a",
  2213 => x"ff49721e",
  2214 => x"d0ff87de",
  2215 => x"78e0c048",
  2216 => x"4f268efc",
  2217 => x"711e731e",
  2218 => x"4966c84b",
  2219 => x"c14a731e",
  2220 => x"ff49a2e0",
  2221 => x"8efc87d8",
  2222 => x"4f264b26",
  2223 => x"4ad4ff1e",
  2224 => x"ff7affc3",
  2225 => x"e1c048d0",
  2226 => x"c47ade78",
  2227 => x"7abfd4d0",
  2228 => x"28c84849",
  2229 => x"48717a70",
  2230 => x"7a7028d0",
  2231 => x"28d84871",
  2232 => x"d0ff7a70",
  2233 => x"78e0c048",
  2234 => x"5e0e4f26",
  2235 => x"0e5d5c5b",
  2236 => x"d0c44c71",
  2237 => x"494dbfd4",
  2238 => x"4b712974",
  2239 => x"c19b66d0",
  2240 => x"b766d483",
  2241 => x"87c204ab",
  2242 => x"66d04bc0",
  2243 => x"ff317449",
  2244 => x"739975b9",
  2245 => x"7232744a",
  2246 => x"c4b07148",
  2247 => x"fe58d8d0",
  2248 => x"4d2687da",
  2249 => x"4b264c26",
  2250 => x"ff1e4f26",
  2251 => x"c9c848d0",
  2252 => x"ff487178",
  2253 => x"267808d4",
  2254 => x"4a711e4f",
  2255 => x"ff87eb49",
  2256 => x"78c848d0",
  2257 => x"731e4f26",
  2258 => x"c44b711e",
  2259 => x"02bfe4d0",
  2260 => x"ebc287c3",
  2261 => x"48d0ff87",
  2262 => x"7378c9c8",
  2263 => x"b1e0c049",
  2264 => x"7148d4ff",
  2265 => x"d8d0c478",
  2266 => x"c878c048",
  2267 => x"87c50266",
  2268 => x"c249ffc3",
  2269 => x"c449c087",
  2270 => x"cc59e0d0",
  2271 => x"87c60266",
  2272 => x"4ad5d5c5",
  2273 => x"ffcf87c4",
  2274 => x"d0c44aff",
  2275 => x"d0c45ae4",
  2276 => x"78c148e4",
  2277 => x"4f264b26",
  2278 => x"5c5b5e0e",
  2279 => x"4d710e5d",
  2280 => x"bfe0d0c4",
  2281 => x"029d754b",
  2282 => x"c84987cb",
  2283 => x"fcccc291",
  2284 => x"c482714a",
  2285 => x"fcd0c287",
  2286 => x"124cc04a",
  2287 => x"c4997349",
  2288 => x"b9bfdcd0",
  2289 => x"7148d4ff",
  2290 => x"2bb7c178",
  2291 => x"acb7c884",
  2292 => x"c487e804",
  2293 => x"48bfd8d0",
  2294 => x"d0c480c8",
  2295 => x"4d2658dc",
  2296 => x"4b264c26",
  2297 => x"731e4f26",
  2298 => x"134b711e",
  2299 => x"cb029a4a",
  2300 => x"fe497287",
  2301 => x"4a1387e2",
  2302 => x"87f5059a",
  2303 => x"4f264b26",
  2304 => x"d8d0c41e",
  2305 => x"d0c449bf",
  2306 => x"a1c148d8",
  2307 => x"b7c0c478",
  2308 => x"87db03a9",
  2309 => x"c448d4ff",
  2310 => x"78bfdcd0",
  2311 => x"bfd8d0c4",
  2312 => x"d8d0c449",
  2313 => x"78a1c148",
  2314 => x"a9b7c0c4",
  2315 => x"ff87e504",
  2316 => x"78c848d0",
  2317 => x"48e4d0c4",
  2318 => x"4f2678c0",
  2319 => x"00000000",
  2320 => x"00000000",
  2321 => x"5f000000",
  2322 => x"0000005f",
  2323 => x"00030300",
  2324 => x"00000303",
  2325 => x"147f7f14",
  2326 => x"00147f7f",
  2327 => x"6b2e2400",
  2328 => x"00123a6b",
  2329 => x"18366a4c",
  2330 => x"0032566c",
  2331 => x"594f7e30",
  2332 => x"40683a77",
  2333 => x"07040000",
  2334 => x"00000003",
  2335 => x"3e1c0000",
  2336 => x"00004163",
  2337 => x"63410000",
  2338 => x"00001c3e",
  2339 => x"1c3e2a08",
  2340 => x"082a3e1c",
  2341 => x"3e080800",
  2342 => x"0008083e",
  2343 => x"e0800000",
  2344 => x"00000060",
  2345 => x"08080800",
  2346 => x"00080808",
  2347 => x"60000000",
  2348 => x"00000060",
  2349 => x"18306040",
  2350 => x"0103060c",
  2351 => x"597f3e00",
  2352 => x"003e7f4d",
  2353 => x"7f060400",
  2354 => x"0000007f",
  2355 => x"71634200",
  2356 => x"00464f59",
  2357 => x"49632200",
  2358 => x"00367f49",
  2359 => x"13161c18",
  2360 => x"00107f7f",
  2361 => x"45672700",
  2362 => x"00397d45",
  2363 => x"4b7e3c00",
  2364 => x"00307949",
  2365 => x"71010100",
  2366 => x"00070f79",
  2367 => x"497f3600",
  2368 => x"00367f49",
  2369 => x"494f0600",
  2370 => x"001e3f69",
  2371 => x"66000000",
  2372 => x"00000066",
  2373 => x"e6800000",
  2374 => x"00000066",
  2375 => x"14080800",
  2376 => x"00222214",
  2377 => x"14141400",
  2378 => x"00141414",
  2379 => x"14222200",
  2380 => x"00080814",
  2381 => x"51030200",
  2382 => x"00060f59",
  2383 => x"5d417f3e",
  2384 => x"001e1f55",
  2385 => x"097f7e00",
  2386 => x"007e7f09",
  2387 => x"497f7f00",
  2388 => x"00367f49",
  2389 => x"633e1c00",
  2390 => x"00414141",
  2391 => x"417f7f00",
  2392 => x"001c3e63",
  2393 => x"497f7f00",
  2394 => x"00414149",
  2395 => x"097f7f00",
  2396 => x"00010109",
  2397 => x"417f3e00",
  2398 => x"007a7b49",
  2399 => x"087f7f00",
  2400 => x"007f7f08",
  2401 => x"7f410000",
  2402 => x"0000417f",
  2403 => x"40602000",
  2404 => x"003f7f40",
  2405 => x"1c087f7f",
  2406 => x"00416336",
  2407 => x"407f7f00",
  2408 => x"00404040",
  2409 => x"0c067f7f",
  2410 => x"007f7f06",
  2411 => x"0c067f7f",
  2412 => x"007f7f18",
  2413 => x"417f3e00",
  2414 => x"003e7f41",
  2415 => x"097f7f00",
  2416 => x"00060f09",
  2417 => x"61417f3e",
  2418 => x"00407e7f",
  2419 => x"097f7f00",
  2420 => x"00667f19",
  2421 => x"4d6f2600",
  2422 => x"00327b59",
  2423 => x"7f010100",
  2424 => x"0001017f",
  2425 => x"407f3f00",
  2426 => x"003f7f40",
  2427 => x"703f0f00",
  2428 => x"000f3f70",
  2429 => x"18307f7f",
  2430 => x"007f7f30",
  2431 => x"1c366341",
  2432 => x"4163361c",
  2433 => x"7c060301",
  2434 => x"0103067c",
  2435 => x"4d597161",
  2436 => x"00414347",
  2437 => x"7f7f0000",
  2438 => x"00004141",
  2439 => x"0c060301",
  2440 => x"40603018",
  2441 => x"41410000",
  2442 => x"00007f7f",
  2443 => x"03060c08",
  2444 => x"00080c06",
  2445 => x"80808080",
  2446 => x"00808080",
  2447 => x"03000000",
  2448 => x"00000407",
  2449 => x"54742000",
  2450 => x"00787c54",
  2451 => x"447f7f00",
  2452 => x"00387c44",
  2453 => x"447c3800",
  2454 => x"00004444",
  2455 => x"447c3800",
  2456 => x"007f7f44",
  2457 => x"547c3800",
  2458 => x"00185c54",
  2459 => x"7f7e0400",
  2460 => x"00000505",
  2461 => x"a4bc1800",
  2462 => x"007cfca4",
  2463 => x"047f7f00",
  2464 => x"00787c04",
  2465 => x"3d000000",
  2466 => x"0000407d",
  2467 => x"80808000",
  2468 => x"00007dfd",
  2469 => x"107f7f00",
  2470 => x"00446c38",
  2471 => x"3f000000",
  2472 => x"0000407f",
  2473 => x"180c7c7c",
  2474 => x"00787c0c",
  2475 => x"047c7c00",
  2476 => x"00787c04",
  2477 => x"447c3800",
  2478 => x"00387c44",
  2479 => x"24fcfc00",
  2480 => x"00183c24",
  2481 => x"243c1800",
  2482 => x"00fcfc24",
  2483 => x"047c7c00",
  2484 => x"00080c04",
  2485 => x"545c4800",
  2486 => x"00207454",
  2487 => x"7f3f0400",
  2488 => x"00004444",
  2489 => x"407c3c00",
  2490 => x"007c7c40",
  2491 => x"603c1c00",
  2492 => x"001c3c60",
  2493 => x"30607c3c",
  2494 => x"003c7c60",
  2495 => x"10386c44",
  2496 => x"00446c38",
  2497 => x"e0bc1c00",
  2498 => x"001c3c60",
  2499 => x"74644400",
  2500 => x"00444c5c",
  2501 => x"3e080800",
  2502 => x"00414177",
  2503 => x"7f000000",
  2504 => x"0000007f",
  2505 => x"77414100",
  2506 => x"0008083e",
  2507 => x"03010102",
  2508 => x"00010202",
  2509 => x"7f7f7f7f",
  2510 => x"007f7f7f",
  2511 => x"1c1c0808",
  2512 => x"7f7f3e3e",
  2513 => x"3e3e7f7f",
  2514 => x"08081c1c",
  2515 => x"7c181000",
  2516 => x"0010187c",
  2517 => x"7c301000",
  2518 => x"0010307c",
  2519 => x"60603010",
  2520 => x"00061e78",
  2521 => x"183c6642",
  2522 => x"0042663c",
  2523 => x"c26a3878",
  2524 => x"00386cc6",
  2525 => x"60000060",
  2526 => x"00600000",
  2527 => x"5c5b5e0e",
  2528 => x"86fc0e5d",
  2529 => x"d0c47e71",
  2530 => x"c04cbff8",
  2531 => x"c41ec04b",
  2532 => x"c402ab66",
  2533 => x"c24dc087",
  2534 => x"754dc187",
  2535 => x"ee49731e",
  2536 => x"86c887e4",
  2537 => x"ef49e0c0",
  2538 => x"a4c487ee",
  2539 => x"f0496a4a",
  2540 => x"cbf187f4",
  2541 => x"c184cc87",
  2542 => x"abb7c883",
  2543 => x"87cdff04",
  2544 => x"4d268efc",
  2545 => x"4b264c26",
  2546 => x"711e4f26",
  2547 => x"fcd0c44a",
  2548 => x"fcd0c45a",
  2549 => x"4978c748",
  2550 => x"2687e1fe",
  2551 => x"1e731e4f",
  2552 => x"b7c04a71",
  2553 => x"87d303aa",
  2554 => x"bfe0eec2",
  2555 => x"c187c405",
  2556 => x"c087c24b",
  2557 => x"e4eec24b",
  2558 => x"c287c45b",
  2559 => x"c25ae4ee",
  2560 => x"4abfe0ee",
  2561 => x"c0c19ac1",
  2562 => x"ecec49a2",
  2563 => x"c248fc87",
  2564 => x"78bfe0ee",
  2565 => x"4f264b26",
  2566 => x"c44a711e",
  2567 => x"49721e66",
  2568 => x"fc87c1ea",
  2569 => x"1e4f268e",
  2570 => x"bfe0eec2",
  2571 => x"cbdfff49",
  2572 => x"f0d0c487",
  2573 => x"78bfe848",
  2574 => x"48ecd0c4",
  2575 => x"c478bfec",
  2576 => x"4abff0d0",
  2577 => x"99ffc349",
  2578 => x"722ab7c8",
  2579 => x"c4b07148",
  2580 => x"2658f8d0",
  2581 => x"5b5e0e4f",
  2582 => x"710e5d5c",
  2583 => x"87c7ff4b",
  2584 => x"48e8d0c4",
  2585 => x"497350c0",
  2586 => x"87f0deff",
  2587 => x"c24c4970",
  2588 => x"49eecb9c",
  2589 => x"87d8d9c1",
  2590 => x"c44d4970",
  2591 => x"bf97e8d0",
  2592 => x"87e5c105",
  2593 => x"c44966d0",
  2594 => x"99bff4d0",
  2595 => x"d487d705",
  2596 => x"d0c44966",
  2597 => x"0599bfec",
  2598 => x"497387cc",
  2599 => x"87fcddff",
  2600 => x"c1029870",
  2601 => x"4cc187c3",
  2602 => x"7587fcfd",
  2603 => x"ebd8c149",
  2604 => x"02987087",
  2605 => x"d0c487c6",
  2606 => x"50c148e8",
  2607 => x"97e8d0c4",
  2608 => x"e4c005bf",
  2609 => x"f4d0c487",
  2610 => x"66d049bf",
  2611 => x"d5ff0599",
  2612 => x"ecd0c487",
  2613 => x"66d449bf",
  2614 => x"c9ff0599",
  2615 => x"ff497387",
  2616 => x"7087f9dc",
  2617 => x"fdfe0598",
  2618 => x"26487487",
  2619 => x"264c264d",
  2620 => x"0e4f264b",
  2621 => x"5d5c5b5e",
  2622 => x"c886f00e",
  2623 => x"78c048a6",
  2624 => x"78c080c4",
  2625 => x"f87ebfec",
  2626 => x"f8d0c480",
  2627 => x"1ec178bf",
  2628 => x"49c71ec0",
  2629 => x"c887fefc",
  2630 => x"02987086",
  2631 => x"49ff87d1",
  2632 => x"c187fafa",
  2633 => x"dbff49da",
  2634 => x"a6c887f2",
  2635 => x"c478c148",
  2636 => x"bf97e8d0",
  2637 => x"c187c402",
  2638 => x"c487fad6",
  2639 => x"4bbff0d0",
  2640 => x"bfe0eec2",
  2641 => x"87c7c105",
  2642 => x"4dc0c0c8",
  2643 => x"4ce4fdc3",
  2644 => x"dbff4914",
  2645 => x"987087c6",
  2646 => x"7587c202",
  2647 => x"2db7c1b3",
  2648 => x"87ecff05",
  2649 => x"ff49fdc3",
  2650 => x"c387f1da",
  2651 => x"daff49fa",
  2652 => x"497387ea",
  2653 => x"7199ffc3",
  2654 => x"fa49c01e",
  2655 => x"497387da",
  2656 => x"7129b7c8",
  2657 => x"fa49c11e",
  2658 => x"86c887ce",
  2659 => x"c487e9c6",
  2660 => x"4bbff4d0",
  2661 => x"e0c0029b",
  2662 => x"dceec287",
  2663 => x"d4c149bf",
  2664 => x"987087fa",
  2665 => x"c087c405",
  2666 => x"c287d44b",
  2667 => x"d4c149e0",
  2668 => x"eec287de",
  2669 => x"c6c058e0",
  2670 => x"dceec287",
  2671 => x"7378c048",
  2672 => x"0599c249",
  2673 => x"ebc387cf",
  2674 => x"cfd9ff49",
  2675 => x"c2497087",
  2676 => x"c5c00299",
  2677 => x"48a6cc87",
  2678 => x"497378fb",
  2679 => x"cf0599c1",
  2680 => x"49f4c387",
  2681 => x"87f4d8ff",
  2682 => x"99c24970",
  2683 => x"87c5c002",
  2684 => x"fa48a6cc",
  2685 => x"c8497378",
  2686 => x"cec00599",
  2687 => x"49f5c387",
  2688 => x"87d8d8ff",
  2689 => x"99c24970",
  2690 => x"c487dc02",
  2691 => x"02bffcd0",
  2692 => x"4887cac0",
  2693 => x"d1c488c1",
  2694 => x"c5c058c0",
  2695 => x"48a6cc87",
  2696 => x"a6c878ff",
  2697 => x"7378c148",
  2698 => x"0599c449",
  2699 => x"c387cfc0",
  2700 => x"d7ff49f2",
  2701 => x"497087e6",
  2702 => x"c00299c2",
  2703 => x"d0c487e2",
  2704 => x"487ebffc",
  2705 => x"03a8b7c7",
  2706 => x"6e87cbc0",
  2707 => x"c480c148",
  2708 => x"c058c0d1",
  2709 => x"a6cc87c5",
  2710 => x"c878fe48",
  2711 => x"78c148a6",
  2712 => x"ff49fdc3",
  2713 => x"7087f5d6",
  2714 => x"0299c249",
  2715 => x"c487dbc0",
  2716 => x"02bffcd0",
  2717 => x"c487c9c0",
  2718 => x"c048fcd0",
  2719 => x"87c5c078",
  2720 => x"fd48a6cc",
  2721 => x"48a6c878",
  2722 => x"fac378c1",
  2723 => x"cbd6ff49",
  2724 => x"c2497087",
  2725 => x"dfc00299",
  2726 => x"fcd0c487",
  2727 => x"b7c748bf",
  2728 => x"c9c003a8",
  2729 => x"fcd0c487",
  2730 => x"c078c748",
  2731 => x"a6cc87c5",
  2732 => x"c878fc48",
  2733 => x"78c148a6",
  2734 => x"c04866cc",
  2735 => x"c003a8b7",
  2736 => x"66c487d6",
  2737 => x"80e0c148",
  2738 => x"bf6e7e70",
  2739 => x"87c8c002",
  2740 => x"cc4bbf6e",
  2741 => x"0f734966",
  2742 => x"f0c31ec0",
  2743 => x"49dac11e",
  2744 => x"c887f2f5",
  2745 => x"02987086",
  2746 => x"c487d9c0",
  2747 => x"7ebffcd0",
  2748 => x"91cc496e",
  2749 => x"714a66c4",
  2750 => x"c0026a82",
  2751 => x"4b6a87c6",
  2752 => x"0f73496e",
  2753 => x"c00266c8",
  2754 => x"d0c487c8",
  2755 => x"f149bffc",
  2756 => x"eec287ea",
  2757 => x"c002bfe4",
  2758 => x"c14987de",
  2759 => x"7087fdce",
  2760 => x"d3c00298",
  2761 => x"fcd0c487",
  2762 => x"cff149bf",
  2763 => x"f249c087",
  2764 => x"eec287eb",
  2765 => x"78c048e4",
  2766 => x"4d268ef0",
  2767 => x"4b264c26",
  2768 => x"5e0e4f26",
  2769 => x"0e5d5c5b",
  2770 => x"4c7186fc",
  2771 => x"bff8d0c4",
  2772 => x"a1d4c149",
  2773 => x"81d8c14d",
  2774 => x"9c747e69",
  2775 => x"c487cf02",
  2776 => x"7b744ba5",
  2777 => x"bff8d0c4",
  2778 => x"87def149",
  2779 => x"9c747b6e",
  2780 => x"c087c405",
  2781 => x"c187c24b",
  2782 => x"f149734b",
  2783 => x"66d487df",
  2784 => x"4987c902",
  2785 => x"87c8cdc1",
  2786 => x"87c24a70",
  2787 => x"eec24ac0",
  2788 => x"8efc5ae8",
  2789 => x"4c264d26",
  2790 => x"4f264b26",
  2791 => x"00000000",
  2792 => x"00000000",
  2793 => x"00000000",
  2794 => x"711e731e",
  2795 => x"cbc1494b",
  2796 => x"d1dafd4a",
  2797 => x"1e4a7087",
  2798 => x"fcc04972",
  2799 => x"c5dafd4a",
  2800 => x"26497087",
  2801 => x"4866c84a",
  2802 => x"49725071",
  2803 => x"fd4afcc0",
  2804 => x"7187f3d9",
  2805 => x"4966c84a",
  2806 => x"517281c1",
  2807 => x"cbc14973",
  2808 => x"e1d9fd4a",
  2809 => x"c84a7187",
  2810 => x"81c24966",
  2811 => x"4b265172",
  2812 => x"731e4f26",
  2813 => x"c84b711e",
  2814 => x"cbc14966",
  2815 => x"4a66cc91",
  2816 => x"4a7349a1",
  2817 => x"92d4c6c1",
  2818 => x"c249a172",
  2819 => x"487189d6",
  2820 => x"4f264b26",
  2821 => x"5c5b5e0e",
  2822 => x"86fc0e5d",
  2823 => x"6b974b71",
  2824 => x"87e4c002",
  2825 => x"487e6b97",
  2826 => x"a8b7f0c0",
  2827 => x"6e87d904",
  2828 => x"b7f9c048",
  2829 => x"87d001a8",
  2830 => x"496e83c1",
  2831 => x"ca89f0c0",
  2832 => x"4866d491",
  2833 => x"87c55071",
  2834 => x"ebc448c0",
  2835 => x"026b9787",
  2836 => x"9787e9c0",
  2837 => x"c0487e6b",
  2838 => x"04a8b7f0",
  2839 => x"486e87de",
  2840 => x"a8b7f9c0",
  2841 => x"c187d501",
  2842 => x"c0496e83",
  2843 => x"66d489f0",
  2844 => x"a14abf97",
  2845 => x"4866d449",
  2846 => x"87c55071",
  2847 => x"f7c348c0",
  2848 => x"026b9787",
  2849 => x"6b9787cd",
  2850 => x"a9fac049",
  2851 => x"c187c405",
  2852 => x"c087c583",
  2853 => x"87e0c348",
  2854 => x"c0026b97",
  2855 => x"6b9787e7",
  2856 => x"f0c0487e",
  2857 => x"dc04a8b7",
  2858 => x"c0486e87",
  2859 => x"01a8b7f9",
  2860 => x"83c187d3",
  2861 => x"f0c0496e",
  2862 => x"d491ca89",
  2863 => x"84c14c66",
  2864 => x"c57c9771",
  2865 => x"c248c087",
  2866 => x"6b9787ee",
  2867 => x"87e4c002",
  2868 => x"487e6b97",
  2869 => x"a8b7f0c0",
  2870 => x"6e87d904",
  2871 => x"b7f9c048",
  2872 => x"87d001a8",
  2873 => x"496e83c1",
  2874 => x"9789f0c0",
  2875 => x"49a14a6c",
  2876 => x"87c57c97",
  2877 => x"ffc148c0",
  2878 => x"026b9787",
  2879 => x"6b9787cd",
  2880 => x"a9fac049",
  2881 => x"c187c405",
  2882 => x"c087c583",
  2883 => x"87e8c148",
  2884 => x"c0026b97",
  2885 => x"6b9787e4",
  2886 => x"b7f0c04a",
  2887 => x"87da04aa",
  2888 => x"aab7f9c0",
  2889 => x"c187d301",
  2890 => x"c0497283",
  2891 => x"91ca89f0",
  2892 => x"c24d66d4",
  2893 => x"7d977185",
  2894 => x"48c087c5",
  2895 => x"9787f9c0",
  2896 => x"e4c0026b",
  2897 => x"7e6b9787",
  2898 => x"b7f0c048",
  2899 => x"87d904a8",
  2900 => x"f9c0486e",
  2901 => x"d001a8b7",
  2902 => x"6e83c187",
  2903 => x"89f0c049",
  2904 => x"a14a6d97",
  2905 => x"c47d9749",
  2906 => x"cb48c087",
  2907 => x"026b9787",
  2908 => x"48c087c4",
  2909 => x"48c187c2",
  2910 => x"4d268efc",
  2911 => x"4b264c26",
  2912 => x"5e0e4f26",
  2913 => x"0e5d5c5b",
  2914 => x"4d7186f8",
  2915 => x"c44b4cc0",
  2916 => x"fd49f8d1",
  2917 => x"7087ccfc",
  2918 => x"aab7c04a",
  2919 => x"87f2c204",
  2920 => x"c202aaca",
  2921 => x"e0c087ec",
  2922 => x"87cf02aa",
  2923 => x"ca02aac9",
  2924 => x"02aacd87",
  2925 => x"aaca87c5",
  2926 => x"7487c605",
  2927 => x"d1c2029c",
  2928 => x"aae2c087",
  2929 => x"7487cc05",
  2930 => x"71b9c149",
  2931 => x"9cffc34c",
  2932 => x"7487fcfe",
  2933 => x"e7c1059c",
  2934 => x"b7e1c187",
  2935 => x"87c804aa",
  2936 => x"aab7fac1",
  2937 => x"87d8c106",
  2938 => x"aab7c1c1",
  2939 => x"c187c804",
  2940 => x"06aab7da",
  2941 => x"c087c9c1",
  2942 => x"04aab7f0",
  2943 => x"f9c087c8",
  2944 => x"c006aab7",
  2945 => x"dbc187fa",
  2946 => x"f3c002aa",
  2947 => x"aaddc187",
  2948 => x"87ecc002",
  2949 => x"02aaedc0",
  2950 => x"c187e5c0",
  2951 => x"df02aadf",
  2952 => x"aaecc087",
  2953 => x"c087d902",
  2954 => x"d302aafd",
  2955 => x"aafec187",
  2956 => x"c087cd02",
  2957 => x"c702aafa",
  2958 => x"aaefc087",
  2959 => x"87cffd05",
  2960 => x"abb7ffc0",
  2961 => x"87c7fd03",
  2962 => x"c149a375",
  2963 => x"fc517283",
  2964 => x"a37587fd",
  2965 => x"b751c049",
  2966 => x"87c403aa",
  2967 => x"87df7ec4",
  2968 => x"c7059b73",
  2969 => x"48a6c487",
  2970 => x"87d078c3",
  2971 => x"c4029c74",
  2972 => x"c27ec187",
  2973 => x"c47ec087",
  2974 => x"786e48a6",
  2975 => x"6e7e66c4",
  2976 => x"268ef848",
  2977 => x"264c264d",
  2978 => x"0e4f264b",
  2979 => x"5d5c5b5e",
  2980 => x"c44d710e",
  2981 => x"c04bc0d1",
  2982 => x"49f8c04a",
  2983 => x"87e9c8fd",
  2984 => x"d1c41e75",
  2985 => x"ebfd49f8",
  2986 => x"86c487dd",
  2987 => x"c5059870",
  2988 => x"c04cc187",
  2989 => x"49c187eb",
  2990 => x"7087f0c0",
  2991 => x"ca059c4c",
  2992 => x"c4d1c487",
  2993 => x"e2c049bf",
  2994 => x"744c7087",
  2995 => x"87cb059c",
  2996 => x"48c0d1c4",
  2997 => x"bfd4d1c4",
  2998 => x"c487c678",
  2999 => x"c048c4d1",
  3000 => x"26487478",
  3001 => x"264c264d",
  3002 => x"0e4f264b",
  3003 => x"5d5c5b5e",
  3004 => x"86ccff0e",
  3005 => x"59a6ecc0",
  3006 => x"974c4dc0",
  3007 => x"48a6c17e",
  3008 => x"80c050c0",
  3009 => x"c080c150",
  3010 => x"c080c478",
  3011 => x"c080c478",
  3012 => x"c080c478",
  3013 => x"c080c478",
  3014 => x"c0d2c478",
  3015 => x"87c505bf",
  3016 => x"d3d048c1",
  3017 => x"f8d1c487",
  3018 => x"d078c048",
  3019 => x"f478c080",
  3020 => x"c4d2c480",
  3021 => x"d0c378bf",
  3022 => x"78c048c0",
  3023 => x"48d4d1c4",
  3024 => x"cfc378c0",
  3025 => x"f9f849c0",
  3026 => x"58a6dc87",
  3027 => x"cd02a8c3",
  3028 => x"4b7587d6",
  3029 => x"87d8029b",
  3030 => x"c1028bc1",
  3031 => x"028b87ee",
  3032 => x"8b87d3c3",
  3033 => x"87f1c602",
  3034 => x"edc7028b",
  3035 => x"87f8cc87",
  3036 => x"cfc34cc0",
  3037 => x"cdc34ac0",
  3038 => x"c3fd49e4",
  3039 => x"987087d1",
  3040 => x"c187c505",
  3041 => x"87e0cc4d",
  3042 => x"4ac0cfc3",
  3043 => x"49eccdc3",
  3044 => x"87fbc2fd",
  3045 => x"c5059870",
  3046 => x"cc4dc287",
  3047 => x"cfc387ca",
  3048 => x"cdc34ac0",
  3049 => x"c2fd49f4",
  3050 => x"987087e5",
  3051 => x"87c5c005",
  3052 => x"f3cb4dc3",
  3053 => x"c0cfc387",
  3054 => x"fccdc34a",
  3055 => x"cec2fd49",
  3056 => x"05987087",
  3057 => x"c487e1cb",
  3058 => x"87dccb4d",
  3059 => x"e0c04874",
  3060 => x"987058a6",
  3061 => x"87cbc105",
  3062 => x"c048a6c8",
  3063 => x"6697c278",
  3064 => x"87cac105",
  3065 => x"bfecd1c4",
  3066 => x"87c7c002",
  3067 => x"50c180fa",
  3068 => x"c387fbc0",
  3069 => x"c41ec0cf",
  3070 => x"fd49e4d1",
  3071 => x"c487c8e6",
  3072 => x"02987086",
  3073 => x"c287c8c0",
  3074 => x"50c148a6",
  3075 => x"c487c3c0",
  3076 => x"fec37e97",
  3077 => x"d1c41eec",
  3078 => x"eafd49f8",
  3079 => x"86c487ef",
  3080 => x"dc87cbc0",
  3081 => x"a8c14866",
  3082 => x"87c2c005",
  3083 => x"84c14dc0",
  3084 => x"c99cffc3",
  3085 => x"a6d487f2",
  3086 => x"66e0c048",
  3087 => x"c0487478",
  3088 => x"7058a6e0",
  3089 => x"fec00598",
  3090 => x"c01eca87",
  3091 => x"c0cfc31e",
  3092 => x"efc4fd49",
  3093 => x"7086c887",
  3094 => x"a6e0c049",
  3095 => x"0266dc59",
  3096 => x"4887d5c0",
  3097 => x"a8b7e3c1",
  3098 => x"87ccc001",
  3099 => x"c14966c4",
  3100 => x"a966dc81",
  3101 => x"87c6c002",
  3102 => x"c27e97c2",
  3103 => x"a6c487d3",
  3104 => x"7866dc48",
  3105 => x"dc87cac2",
  3106 => x"a8c14866",
  3107 => x"87c1c205",
  3108 => x"4ac0cfc3",
  3109 => x"49c4cdc3",
  3110 => x"87f3fefc",
  3111 => x"c0059870",
  3112 => x"e0c087cf",
  3113 => x"e4c048a6",
  3114 => x"80c478f0",
  3115 => x"c5c178c0",
  3116 => x"c0cfc387",
  3117 => x"cccdc34a",
  3118 => x"d2fefc49",
  3119 => x"05987087",
  3120 => x"c087cfc0",
  3121 => x"c048a6e0",
  3122 => x"c478f0e4",
  3123 => x"c078c180",
  3124 => x"cfc387e4",
  3125 => x"cdc34ac0",
  3126 => x"fdfc49d8",
  3127 => x"987087f1",
  3128 => x"87cfc005",
  3129 => x"48a6e0c0",
  3130 => x"78c0e0c0",
  3131 => x"78c180c4",
  3132 => x"c287c3c0",
  3133 => x"e8c07e97",
  3134 => x"66c44866",
  3135 => x"cec005a8",
  3136 => x"dcd1c487",
  3137 => x"66e0c048",
  3138 => x"c080fc78",
  3139 => x"c07866e4",
  3140 => x"c384c14d",
  3141 => x"cfc69cff",
  3142 => x"a6ecc087",
  3143 => x"c0cfc31e",
  3144 => x"87f0eb49",
  3145 => x"987086c4",
  3146 => x"87c6c005",
  3147 => x"c07e97c2",
  3148 => x"eec087e3",
  3149 => x"1e496697",
  3150 => x"6697f1c0",
  3151 => x"f4c01e49",
  3152 => x"ea496697",
  3153 => x"86c887ec",
  3154 => x"d6c24970",
  3155 => x"c8487181",
  3156 => x"a6cc8066",
  3157 => x"c54dc058",
  3158 => x"487487ce",
  3159 => x"58a6e0c0",
  3160 => x"c0059870",
  3161 => x"1eca87d7",
  3162 => x"cfc31ec0",
  3163 => x"c0fd49c0",
  3164 => x"86c887d2",
  3165 => x"a6c54970",
  3166 => x"e6c45997",
  3167 => x"4866dc87",
  3168 => x"c405a8c1",
  3169 => x"ecc087dd",
  3170 => x"cfc31ea6",
  3171 => x"c3ea49c0",
  3172 => x"7086c487",
  3173 => x"c6c00598",
  3174 => x"7e97c287",
  3175 => x"c087c2c4",
  3176 => x"496697ee",
  3177 => x"97f1c01e",
  3178 => x"c01e4966",
  3179 => x"496697f4",
  3180 => x"c887ffe8",
  3181 => x"a6e0c086",
  3182 => x"6697c158",
  3183 => x"a6f4c048",
  3184 => x"05987058",
  3185 => x"c087e7c0",
  3186 => x"c14966e8",
  3187 => x"a966c481",
  3188 => x"87cdc305",
  3189 => x"bfd4d1c4",
  3190 => x"87c5c305",
  3191 => x"c24966dc",
  3192 => x"487181d6",
  3193 => x"c48066c8",
  3194 => x"c258d8d1",
  3195 => x"f0c087f3",
  3196 => x"a8c14866",
  3197 => x"87e9c205",
  3198 => x"c04866c4",
  3199 => x"05a866e8",
  3200 => x"dc87cfc0",
  3201 => x"d6c24966",
  3202 => x"c8487181",
  3203 => x"d1c48066",
  3204 => x"66c458d4",
  3205 => x"a8b7c148",
  3206 => x"87ddc106",
  3207 => x"cc4866dc",
  3208 => x"f4c08866",
  3209 => x"66c458a6",
  3210 => x"66e8c048",
  3211 => x"d0c005a8",
  3212 => x"66f0c087",
  3213 => x"9166d449",
  3214 => x"66d04871",
  3215 => x"d0d1c480",
  3216 => x"66e8c058",
  3217 => x"c481c149",
  3218 => x"c005a966",
  3219 => x"d1c487d9",
  3220 => x"c005bfd4",
  3221 => x"66dc87d1",
  3222 => x"81d6c249",
  3223 => x"718166c8",
  3224 => x"c488c148",
  3225 => x"c058d8d1",
  3226 => x"d44966f0",
  3227 => x"48719166",
  3228 => x"d48066d0",
  3229 => x"e2c058a6",
  3230 => x"4966dc87",
  3231 => x"d481d6c2",
  3232 => x"48719166",
  3233 => x"d48066d0",
  3234 => x"e8c058a6",
  3235 => x"a8c14866",
  3236 => x"87c7c005",
  3237 => x"48ccd1c4",
  3238 => x"cc7866d0",
  3239 => x"66dc48a6",
  3240 => x"c14dc078",
  3241 => x"9cffc384",
  3242 => x"c44866d8",
  3243 => x"c6c002a8",
  3244 => x"026e9787",
  3245 => x"c287cbf2",
  3246 => x"c0056697",
  3247 => x"97c487c6",
  3248 => x"87f6c07e",
  3249 => x"c04866c4",
  3250 => x"05a866e8",
  3251 => x"c487ebc0",
  3252 => x"4abfccd1",
  3253 => x"bfecd1c4",
  3254 => x"70887248",
  3255 => x"dcd1c44a",
  3256 => x"1e7249bf",
  3257 => x"fc4a0972",
  3258 => x"7087e7fc",
  3259 => x"c44a2649",
  3260 => x"48bfd0d1",
  3261 => x"d1c48071",
  3262 => x"66c458d8",
  3263 => x"66e8c048",
  3264 => x"c003a8b7",
  3265 => x"97c487c3",
  3266 => x"026e977e",
  3267 => x"c487c9c0",
  3268 => x"c048c4d1",
  3269 => x"87c7c078",
  3270 => x"48c4d1c4",
  3271 => x"c07866c4",
  3272 => x"c41ea6ec",
  3273 => x"49bfd0d1",
  3274 => x"c487fde1",
  3275 => x"e0d1c486",
  3276 => x"66e8c048",
  3277 => x"486e9778",
  3278 => x"268eccff",
  3279 => x"264c264d",
  3280 => x"004f264b",
  3281 => x"49445541",
  3282 => x"0000004f",
  3283 => x"45444f4d",
  3284 => x"33322f31",
  3285 => x"00003235",
  3286 => x"45444f4d",
  3287 => x"30322f31",
  3288 => x"00003834",
  3289 => x"454c4946",
  3290 => x"00000000",
  3291 => x"43415254",
  3292 => x"0000004b",
  3293 => x"47455250",
  3294 => x"00005041",
  3295 => x"45444e49",
  3296 => x"5e0e0058",
  3297 => x"710e5c5b",
  3298 => x"c44bc14c",
  3299 => x"b7bfd0d1",
  3300 => x"87d004ac",
  3301 => x"bfd4d1c4",
  3302 => x"c701acb7",
  3303 => x"e0d1c487",
  3304 => x"87d348bf",
  3305 => x"c2ed4973",
  3306 => x"c483c187",
  3307 => x"b7bfc4d1",
  3308 => x"d6ff06ab",
  3309 => x"2648ff87",
  3310 => x"264b264c",
  3311 => x"0000004f",
  3312 => x"00000000",
  3313 => x"00000000",
  3314 => x"00000000",
  3315 => x"00000000",
  3316 => x"00000000",
  3317 => x"00000000",
  3318 => x"00000000",
  3319 => x"00000000",
  3320 => x"00000000",
  3321 => x"00000000",
  3322 => x"00000000",
  3323 => x"00000000",
  3324 => x"00000000",
  3325 => x"00000000",
  3326 => x"00000000",
  3327 => x"00000000",
  3328 => x"00000000",
  3329 => x"711e731e",
  3330 => x"721e4a4b",
  3331 => x"fc4aca49",
  3332 => x"7087f3f8",
  3333 => x"d04a2649",
  3334 => x"721e7191",
  3335 => x"fc4aca49",
  3336 => x"7187e3f8",
  3337 => x"7249264a",
  3338 => x"ffc349a1",
  3339 => x"26487199",
  3340 => x"1e4f264b",
  3341 => x"4b711e73",
  3342 => x"b7c4494a",
  3343 => x"cf91ca29",
  3344 => x"49a1729a",
  3345 => x"7199ffc3",
  3346 => x"264b2648",
  3347 => x"1e731e4f",
  3348 => x"ff494a71",
  3349 => x"497087dd",
  3350 => x"c2059b4b",
  3351 => x"c44bc187",
  3352 => x"b7bfc4d1",
  3353 => x"87c106ab",
  3354 => x"e949734b",
  3355 => x"487387fd",
  3356 => x"4f264b26",
  3357 => x"c0f7c41e",
  3358 => x"f6c45997",
  3359 => x"66c448fd",
  3360 => x"5066c850",
  3361 => x"265066cc",
  3362 => x"1e731e4f",
  3363 => x"d0ff4b71",
  3364 => x"78c5c848",
  3365 => x"c148d4ff",
  3366 => x"497378e1",
  3367 => x"2ab7c84a",
  3368 => x"ffc37872",
  3369 => x"ff787199",
  3370 => x"78c448d0",
  3371 => x"4f264b26",
  3372 => x"fef7c41e",
  3373 => x"f7c4599f",
  3374 => x"78c148cc",
  3375 => x"5e0e4f26",
  3376 => x"710e5c5b",
  3377 => x"48d0ff4c",
  3378 => x"ff78c5c8",
  3379 => x"e4c148d4",
  3380 => x"4966cc78",
  3381 => x"9affc34a",
  3382 => x"66cc7872",
  3383 => x"c32ac84a",
  3384 => x"66d09aff",
  3385 => x"7333c74b",
  3386 => x"717872b2",
  3387 => x"fc49741e",
  3388 => x"ff87c4f6",
  3389 => x"78c448d0",
  3390 => x"4c268efc",
  3391 => x"4f264b26",
  3392 => x"c01e731e",
  3393 => x"c44bc0e0",
  3394 => x"02bfd8d1",
  3395 => x"c487e7c1",
  3396 => x"48bfd8f7",
  3397 => x"04a8b7c0",
  3398 => x"c487dbc1",
  3399 => x"abbfdcd1",
  3400 => x"c487d302",
  3401 => x"49bff4d1",
  3402 => x"1e7181d0",
  3403 => x"49e4d1c4",
  3404 => x"87e9d7fd",
  3405 => x"1e7386c4",
  3406 => x"1eccd2c4",
  3407 => x"49e4d1c4",
  3408 => x"87c2d9fd",
  3409 => x"d1c486c8",
  3410 => x"02abbfdc",
  3411 => x"c04987d6",
  3412 => x"c489d0e0",
  3413 => x"81bff4d1",
  3414 => x"d1c41e71",
  3415 => x"d6fd49e4",
  3416 => x"86c487fb",
  3417 => x"1e4966c8",
  3418 => x"d2c41e73",
  3419 => x"cdfd49cc",
  3420 => x"c086c887",
  3421 => x"e4c087e1",
  3422 => x"d2c41ef0",
  3423 => x"d1c41ecc",
  3424 => x"d8fd49e4",
  3425 => x"66d087c0",
  3426 => x"e4c01e49",
  3427 => x"d2c41ef0",
  3428 => x"e9fc49cc",
  3429 => x"2686d087",
  3430 => x"1e4f264b",
  3431 => x"bfecd1c4",
  3432 => x"c487db05",
  3433 => x"c148c4f7",
  3434 => x"1e1ec050",
  3435 => x"49c21ecb",
  3436 => x"cc87c1fb",
  3437 => x"fb49c186",
  3438 => x"48c087cf",
  3439 => x"48c187c2",
  3440 => x"5e0e4f26",
  3441 => x"c00e5c5b",
  3442 => x"c44cf0e4",
  3443 => x"48bfc0f7",
  3444 => x"c006a8c0",
  3445 => x"fbc387e9",
  3446 => x"c049bfcc",
  3447 => x"7087fde3",
  3448 => x"dfc70298",
  3449 => x"c049cd87",
  3450 => x"7087e5e3",
  3451 => x"d0fbc349",
  3452 => x"c0f7c459",
  3453 => x"88c148bf",
  3454 => x"58c4f7c4",
  3455 => x"c487c5c7",
  3456 => x"bf97c4f7",
  3457 => x"05aac24a",
  3458 => x"c487cac3",
  3459 => x"48bfd4f7",
  3460 => x"bfc4d1c4",
  3461 => x"c906a8b7",
  3462 => x"c4f7c487",
  3463 => x"c650c048",
  3464 => x"f7c487e2",
  3465 => x"02bf97d1",
  3466 => x"c487d9c6",
  3467 => x"05bfecd1",
  3468 => x"f7c487da",
  3469 => x"50c148c4",
  3470 => x"cb1e1ec0",
  3471 => x"f849c21e",
  3472 => x"86cc87f2",
  3473 => x"e7f949c1",
  3474 => x"87f8c587",
  3475 => x"48d1f7c4",
  3476 => x"d1c450c0",
  3477 => x"cd02bfd8",
  3478 => x"c01ec187",
  3479 => x"fa49c0e0",
  3480 => x"86c487de",
  3481 => x"f7c487d5",
  3482 => x"c448bfd8",
  3483 => x"b7bfd0d1",
  3484 => x"c6c004a8",
  3485 => x"c5f7c487",
  3486 => x"c450c048",
  3487 => x"48bfdcf7",
  3488 => x"f7c488c1",
  3489 => x"987058e0",
  3490 => x"87cbc005",
  3491 => x"dff849c0",
  3492 => x"c4f7c487",
  3493 => x"c450c048",
  3494 => x"48bfd8f7",
  3495 => x"f7c480c1",
  3496 => x"d1c458dc",
  3497 => x"a8b7bfd4",
  3498 => x"87d8c404",
  3499 => x"bfd4f7c4",
  3500 => x"c480c148",
  3501 => x"7058d8f7",
  3502 => x"87efe049",
  3503 => x"48c5f7c4",
  3504 => x"d1c450c1",
  3505 => x"1e49bfcc",
  3506 => x"49e4d1c4",
  3507 => x"87cdd1fd",
  3508 => x"efc386c4",
  3509 => x"05aac387",
  3510 => x"c487e9c3",
  3511 => x"05bfecd1",
  3512 => x"c487dac0",
  3513 => x"c148c4f7",
  3514 => x"1e1ec050",
  3515 => x"49c21ecb",
  3516 => x"cc87c1f6",
  3517 => x"f649c186",
  3518 => x"c7c387f6",
  3519 => x"d8f7c487",
  3520 => x"fdf149bf",
  3521 => x"d8f7c487",
  3522 => x"d2f7c458",
  3523 => x"c105bf97",
  3524 => x"4bc087d1",
  3525 => x"bff4f7c4",
  3526 => x"a8b7c048",
  3527 => x"87c3c104",
  3528 => x"bfd8d1c4",
  3529 => x"87e4c005",
  3530 => x"bfd8f7c4",
  3531 => x"d0d1c449",
  3532 => x"917489bf",
  3533 => x"bfccd1c4",
  3534 => x"c41e7181",
  3535 => x"fd49e4d1",
  3536 => x"c087dacf",
  3537 => x"f649741e",
  3538 => x"86c887f6",
  3539 => x"bfd8f7c4",
  3540 => x"c480c148",
  3541 => x"c158dcf7",
  3542 => x"f4f7c483",
  3543 => x"06abb7bf",
  3544 => x"c487fdfe",
  3545 => x"c048f4f7",
  3546 => x"d8f7c478",
  3547 => x"f7c448bf",
  3548 => x"a8b7bff0",
  3549 => x"87d7c003",
  3550 => x"bfd8d1c4",
  3551 => x"87cfc005",
  3552 => x"bfd4f7c4",
  3553 => x"c4d1c448",
  3554 => x"06a8b7bf",
  3555 => x"c487f5c0",
  3556 => x"bf97f8f7",
  3557 => x"05a9c149",
  3558 => x"c487d2c0",
  3559 => x"c448d8f7",
  3560 => x"78bfecf7",
  3561 => x"48c0f7c4",
  3562 => x"c6c078c2",
  3563 => x"c4f7c487",
  3564 => x"c450c048",
  3565 => x"bf97f8f7",
  3566 => x"05a9c249",
  3567 => x"c087c5c0",
  3568 => x"87ecf349",
  3569 => x"4b264c26",
  3570 => x"5e0e4f26",
  3571 => x"0e5d5c5b",
  3572 => x"7686c4ff",
  3573 => x"c04ac04b",
  3574 => x"e3fc49e0",
  3575 => x"d0ff87eb",
  3576 => x"78c5c848",
  3577 => x"c148d4ff",
  3578 => x"4dc078e2",
  3579 => x"7cc04c70",
  3580 => x"49a6e0c0",
  3581 => x"516c8175",
  3582 => x"b7cc85c1",
  3583 => x"87ee04ad",
  3584 => x"c448d0ff",
  3585 => x"97e0c078",
  3586 => x"029c4c66",
  3587 => x"c387f3c0",
  3588 => x"fec0028c",
  3589 => x"028cc587",
  3590 => x"cd87e7c6",
  3591 => x"f3c8028c",
  3592 => x"8cc3c387",
  3593 => x"87c5c902",
  3594 => x"cc028cc1",
  3595 => x"028c87e9",
  3596 => x"c387eed0",
  3597 => x"ffd0028c",
  3598 => x"028cc187",
  3599 => x"d487f8c1",
  3600 => x"d6f587f1",
  3601 => x"02987087",
  3602 => x"c087c2d5",
  3603 => x"87f9f049",
  3604 => x"d287fad4",
  3605 => x"a6c17e97",
  3606 => x"50c0c248",
  3607 => x"c150f0c1",
  3608 => x"fcf6c480",
  3609 => x"c450bf97",
  3610 => x"c450ca80",
  3611 => x"fdf6c480",
  3612 => x"c450bf97",
  3613 => x"bf97fef6",
  3614 => x"fff6c450",
  3615 => x"c450bf97",
  3616 => x"c048fff6",
  3617 => x"fef6c450",
  3618 => x"fff6c448",
  3619 => x"c450bf97",
  3620 => x"c448fdf6",
  3621 => x"bf97fef6",
  3622 => x"fcf6c450",
  3623 => x"fdf6c448",
  3624 => x"c150bf97",
  3625 => x"ca1ed21e",
  3626 => x"d1f049a6",
  3627 => x"c086c887",
  3628 => x"87d5ef49",
  3629 => x"f387d6d3",
  3630 => x"987087e1",
  3631 => x"87cdd302",
  3632 => x"6697e1c0",
  3633 => x"a6f0c048",
  3634 => x"02987058",
  3635 => x"c14887da",
  3636 => x"a6f0c088",
  3637 => x"02987058",
  3638 => x"4887edc0",
  3639 => x"f0c088c1",
  3640 => x"987058a6",
  3641 => x"87ecc102",
  3642 => x"c17e97c2",
  3643 => x"c0c248a6",
  3644 => x"c450c150",
  3645 => x"49bfc4d1",
  3646 => x"c387c9ec",
  3647 => x"c05008a6",
  3648 => x"c248a6ec",
  3649 => x"87e4c278",
  3650 => x"bfc0d1c4",
  3651 => x"81d6c249",
  3652 => x"1ea6f0c0",
  3653 => x"cfcaff71",
  3654 => x"9786c487",
  3655 => x"48a6c17e",
  3656 => x"c050c0c2",
  3657 => x"496697f0",
  3658 => x"c287d9eb",
  3659 => x"c05008a6",
  3660 => x"496697f1",
  3661 => x"c387cdeb",
  3662 => x"c05008a6",
  3663 => x"496697f2",
  3664 => x"c487c1eb",
  3665 => x"c55008a6",
  3666 => x"50c048a6",
  3667 => x"c480e6c0",
  3668 => x"87d8c178",
  3669 => x"6697e2c0",
  3670 => x"87f1eb49",
  3671 => x"bfd0d1c4",
  3672 => x"81d6c249",
  3673 => x"1ea6f0c0",
  3674 => x"fbc8ff71",
  3675 => x"9786c487",
  3676 => x"48a6c17e",
  3677 => x"c050c0c2",
  3678 => x"496697f0",
  3679 => x"c287c5ea",
  3680 => x"c05008a6",
  3681 => x"496697f1",
  3682 => x"c387f9e9",
  3683 => x"c05008a6",
  3684 => x"496697f2",
  3685 => x"c487ede9",
  3686 => x"c45008a6",
  3687 => x"49bfd8d1",
  3688 => x"a6c931c2",
  3689 => x"c0485997",
  3690 => x"78c480e7",
  3691 => x"f0c01ec1",
  3692 => x"a6ca1e66",
  3693 => x"87c6ec49",
  3694 => x"49c086c8",
  3695 => x"cf87caeb",
  3696 => x"d6ef87cb",
  3697 => x"02987087",
  3698 => x"c087c2cf",
  3699 => x"496697e1",
  3700 => x"e2c031d0",
  3701 => x"c84a6697",
  3702 => x"c0b17232",
  3703 => x"4a6697e3",
  3704 => x"c74871b1",
  3705 => x"98ffffff",
  3706 => x"58a6f0c0",
  3707 => x"6697e4c0",
  3708 => x"87c8c002",
  3709 => x"a6f8c048",
  3710 => x"87c7c058",
  3711 => x"48a6f4c0",
  3712 => x"c078c0c4",
  3713 => x"e54966ec",
  3714 => x"f7c487f8",
  3715 => x"f7c458d8",
  3716 => x"78c048c0",
  3717 => x"48d8f7c4",
  3718 => x"4066ecc0",
  3719 => x"7866f4c0",
  3720 => x"4966ecc0",
  3721 => x"bfd0d1c4",
  3722 => x"dcd1c489",
  3723 => x"d1c491bf",
  3724 => x"7181bfcc",
  3725 => x"e4d1c41e",
  3726 => x"e0c3fd49",
  3727 => x"c486c487",
  3728 => x"c048e8f7",
  3729 => x"d1f7c478",
  3730 => x"c450c148",
  3731 => x"c248c4f7",
  3732 => x"87f9cc50",
  3733 => x"6697e4c0",
  3734 => x"87c9c002",
  3735 => x"48d0f7c4",
  3736 => x"e8cc50c1",
  3737 => x"e849c087",
  3738 => x"e0cc87df",
  3739 => x"87ebec87",
  3740 => x"cc029870",
  3741 => x"e9c087d7",
  3742 => x"48496697",
  3743 => x"c098c0c3",
  3744 => x"7058a6f0",
  3745 => x"dcc00298",
  3746 => x"c0c14887",
  3747 => x"a6f0c088",
  3748 => x"02987058",
  3749 => x"4887edc0",
  3750 => x"c088c0c1",
  3751 => x"7058a6f0",
  3752 => x"cdc10298",
  3753 => x"97e3c087",
  3754 => x"31d04966",
  3755 => x"6697e4c0",
  3756 => x"7232c84a",
  3757 => x"97e5c0b1",
  3758 => x"71484a66",
  3759 => x"a6f0c0b0",
  3760 => x"87ffc058",
  3761 => x"6697e4c0",
  3762 => x"87e7e549",
  3763 => x"c01e4970",
  3764 => x"496697e7",
  3765 => x"7087dce5",
  3766 => x"eac01e49",
  3767 => x"e5496697",
  3768 => x"4a7087d1",
  3769 => x"c9c4ff49",
  3770 => x"c086c887",
  3771 => x"c058a6f0",
  3772 => x"e2c087d1",
  3773 => x"e5496697",
  3774 => x"ecc087d3",
  3775 => x"d1c448a6",
  3776 => x"c478bfd0",
  3777 => x"c048c0f7",
  3778 => x"d8f7c478",
  3779 => x"66ecc048",
  3780 => x"ede14978",
  3781 => x"d8f7c487",
  3782 => x"ecf7c458",
  3783 => x"66ecc048",
  3784 => x"c0d1c440",
  3785 => x"f7c478bf",
  3786 => x"e1c048f8",
  3787 => x"c4506697",
  3788 => x"c148f4f7",
  3789 => x"f8f7c478",
  3790 => x"9949bf97",
  3791 => x"87c9c005",
  3792 => x"48c4f7c4",
  3793 => x"c6c050c4",
  3794 => x"c4f7c487",
  3795 => x"c050c348",
  3796 => x"87dce549",
  3797 => x"e987f6c8",
  3798 => x"987087c1",
  3799 => x"87edc802",
  3800 => x"6697e9c0",
  3801 => x"c0c34849",
  3802 => x"a6f0c098",
  3803 => x"02987058",
  3804 => x"4887dcc0",
  3805 => x"c088c0c1",
  3806 => x"7058a6f0",
  3807 => x"edc00298",
  3808 => x"c0c14887",
  3809 => x"a6f0c088",
  3810 => x"02987058",
  3811 => x"c087cdc1",
  3812 => x"496697e3",
  3813 => x"e4c031d0",
  3814 => x"c84a6697",
  3815 => x"c0b17232",
  3816 => x"4a6697e5",
  3817 => x"c0b07148",
  3818 => x"c158a6f0",
  3819 => x"e4c087f4",
  3820 => x"e1496697",
  3821 => x"497087fd",
  3822 => x"97e7c01e",
  3823 => x"f2e14966",
  3824 => x"1e497087",
  3825 => x"6697eac0",
  3826 => x"87e7e149",
  3827 => x"ff494a70",
  3828 => x"c887dfc0",
  3829 => x"a6f0c086",
  3830 => x"87c6c158",
  3831 => x"6697e2c0",
  3832 => x"87cfe149",
  3833 => x"c0484970",
  3834 => x"7058a6f0",
  3835 => x"c6c00598",
  3836 => x"a6ecc087",
  3837 => x"c078c148",
  3838 => x"c44866ec",
  3839 => x"b7bfc4d1",
  3840 => x"ccc006a8",
  3841 => x"a6f4c087",
  3842 => x"c0d1c448",
  3843 => x"c9c078bf",
  3844 => x"a6f4c087",
  3845 => x"d4d1c448",
  3846 => x"ecc078bf",
  3847 => x"f4c048a6",
  3848 => x"f7c47866",
  3849 => x"e1c048f8",
  3850 => x"c4506697",
  3851 => x"c048f0f7",
  3852 => x"c47866ec",
  3853 => x"bf97f8f7",
  3854 => x"c0059949",
  3855 => x"f7c487c9",
  3856 => x"50c048c4",
  3857 => x"c487c6c0",
  3858 => x"c348c4f7",
  3859 => x"f8f7c450",
  3860 => x"c249bf97",
  3861 => x"f4c402a9",
  3862 => x"e049c087",
  3863 => x"ecc487eb",
  3864 => x"87f7e487",
  3865 => x"c4029870",
  3866 => x"f7c487e3",
  3867 => x"50c448c4",
  3868 => x"d4e049c0",
  3869 => x"87d5c487",
  3870 => x"7087e0e4",
  3871 => x"ccc40298",
  3872 => x"d8f7c487",
  3873 => x"d1c448bf",
  3874 => x"c088bfd0",
  3875 => x"ca58a6f0",
  3876 => x"a6c17e97",
  3877 => x"50c0c248",
  3878 => x"97c4f7c4",
  3879 => x"f8c048bf",
  3880 => x"a8c458a6",
  3881 => x"87c9c005",
  3882 => x"48a6f4c0",
  3883 => x"e1c078c2",
  3884 => x"66f4c087",
  3885 => x"05a8c348",
  3886 => x"c087c9c0",
  3887 => x"c048a6f8",
  3888 => x"87c6c078",
  3889 => x"48a6f8c0",
  3890 => x"f4c078c3",
  3891 => x"f8c048a6",
  3892 => x"a6c27866",
  3893 => x"66f4c048",
  3894 => x"c450c050",
  3895 => x"49bfd4f7",
  3896 => x"dcff81c1",
  3897 => x"a6c487de",
  3898 => x"f7c45008",
  3899 => x"ff49bfd4",
  3900 => x"c587d1dc",
  3901 => x"c05008a6",
  3902 => x"1e4ba6f0",
  3903 => x"4966f0c0",
  3904 => x"87e4fafe",
  3905 => x"6697f4c0",
  3906 => x"f7dbff49",
  3907 => x"08a6ca87",
  3908 => x"97f5c050",
  3909 => x"dbff4966",
  3910 => x"a6cb87ea",
  3911 => x"f6c05008",
  3912 => x"ff496697",
  3913 => x"cc87dddb",
  3914 => x"735008a6",
  3915 => x"d8f7c41e",
  3916 => x"f9fe49bf",
  3917 => x"f8c087f2",
  3918 => x"ff496697",
  3919 => x"d187c5db",
  3920 => x"c05008a6",
  3921 => x"496697f9",
  3922 => x"87f8daff",
  3923 => x"5008a6d2",
  3924 => x"6697fac0",
  3925 => x"ebdaff49",
  3926 => x"08a6d387",
  3927 => x"ca1ec150",
  3928 => x"49a6d21e",
  3929 => x"87d6ddff",
  3930 => x"49c086d0",
  3931 => x"87d9dcff",
  3932 => x"c087dac0",
  3933 => x"e0c01e1e",
  3934 => x"ff49c51e",
  3935 => x"cc87f5db",
  3936 => x"ccf7c486",
  3937 => x"c178c048",
  3938 => x"fcdbff49",
  3939 => x"8ec4ff87",
  3940 => x"4c264d26",
  3941 => x"4f264b26",
  3942 => x"f41e731e",
  3943 => x"4bd4ff86",
  3944 => x"c848d0ff",
  3945 => x"e3c178c5",
  3946 => x"c04ac07b",
  3947 => x"7249767b",
  3948 => x"c1516b81",
  3949 => x"aab7ca82",
  3950 => x"ff87f004",
  3951 => x"78c448d0",
  3952 => x"4b268ef4",
  3953 => x"c41e4f26",
  3954 => x"c148d1f7",
  3955 => x"1e4f2650",
  3956 => x"48c0f7c4",
  3957 => x"f7c478c0",
  3958 => x"40c048d4",
  3959 => x"e0f7c478",
  3960 => x"c478c048",
  3961 => x"c148c5f7",
  3962 => x"ecd1c450",
  3963 => x"87c402bf",
  3964 => x"87c249c0",
  3965 => x"f7c449c1",
  3966 => x"c45997c8",
  3967 => x"c048e4f7",
  3968 => x"f7c47840",
  3969 => x"40c048cc",
  3970 => x"f7c45050",
  3971 => x"40c048ec",
  3972 => x"f8f7c478",
  3973 => x"c450c048",
  3974 => x"c048faf7",
  3975 => x"f7c4789f",
  3976 => x"50c148d2",
  3977 => x"731e4f26",
  3978 => x"48d0ff1e",
  3979 => x"ff78c5c8",
  3980 => x"e0c148d4",
  3981 => x"c3496878",
  3982 => x"d0ff99ff",
  3983 => x"7178c448",
  3984 => x"99c1494b",
  3985 => x"e687c302",
  3986 => x"497387c0",
  3987 => x"c30299c2",
  3988 => x"87c4fd87",
  3989 => x"99c44973",
  3990 => x"fd87c302",
  3991 => x"497387e8",
  3992 => x"d60299c8",
  3993 => x"87e7fd87",
  3994 => x"c848d0ff",
  3995 => x"d4ff78c5",
  3996 => x"78e6c148",
  3997 => x"d0ff78c0",
  3998 => x"7378c448",
  3999 => x"c499d049",
  4000 => x"5997d6f7",
  4001 => x"87fadcff",
  4002 => x"bfccf7c4",
  4003 => x"c487d702",
  4004 => x"05bfc0f7",
  4005 => x"f7c487d0",
  4006 => x"49bf9ffa",
  4007 => x"87e9d7ff",
  4008 => x"48ccf7c4",
  4009 => x"f7c478c0",
  4010 => x"02bf97d0",
  4011 => x"d0ff87d9",
  4012 => x"78c5c848",
  4013 => x"c148d4ff",
  4014 => x"78c078e5",
  4015 => x"c448d0ff",
  4016 => x"d0f7c478",
  4017 => x"2650c048",
  4018 => x"004f264b",
  4019 => x"00000000",
  4020 => x"ff4a711e",
  4021 => x"7249bfc8",
  4022 => x"4f2648a1",
  4023 => x"bfc8ff1e",
  4024 => x"c0c0fe89",
  4025 => x"a9c0c0c0",
  4026 => x"c087c401",
  4027 => x"c187c24a",
  4028 => x"2648724a",
  4029 => x"fdc31e4f",
  4030 => x"c149bfc4",
  4031 => x"c8fdc3b9",
  4032 => x"48d4ff59",
  4033 => x"ff78ffc3",
  4034 => x"e1c048d0",
  4035 => x"48d4ff78",
  4036 => x"31c478c1",
  4037 => x"d0ff7871",
  4038 => x"78e0c048",
  4039 => x"c31e4f26",
  4040 => x"c41ef8fc",
  4041 => x"fc49e8cb",
  4042 => x"c487dce9",
  4043 => x"02987086",
  4044 => x"c0ff87c3",
  4045 => x"004f2687",
  4046 => x"484b3531",
  4047 => x"2020205a",
  4048 => x"00474643",
  4049 => x"00000000",
  4050 => x"dcf2c11e",
  4051 => x"c150c148",
  4052 => x"c148ccc6",
  4053 => x"f4fdc350",
  4054 => x"c8fd49bf",
  4055 => x"48c087ef",
  4056 => x"00004f26",
  4057 => x"11141258",
  4058 => x"231c1b1d",
  4059 => x"9194595a",
  4060 => x"f4ebf2f5",
  4061 => x"00003f78",
  4062 => x"4f545541",
  4063 => x"544f4f42",
  4064 => x"00584753",
  others => ( x"00000000")
);

-- Xilinx Vivado attributes
attribute ram_style: string;
attribute ram_style of ram: signal is "block";

signal q_local : std_logic_vector((NB_COL * COL_WIDTH)-1 downto 0);

signal wea : std_logic_vector(NB_COL - 1 downto 0);

begin

	output:
	for i in 0 to NB_COL - 1 generate
		q((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= q_local((i+1) * COL_WIDTH - 1 downto i * COL_WIDTH);
	end generate;
    
    -- Generate write enable signals
    -- The Block ram generator doesn't like it when the compare is done in the if statement it self.
    wea <= bytesel when we = '1' else (others => '0');

    process(clk)
    begin
        if rising_edge(clk) then
            q_local <= ram(to_integer(unsigned(addr)));
            for i in 0 to NB_COL - 1 loop
                if (wea(NB_COL-i-1) = '1') then
                    ram(to_integer(unsigned(addr)))((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH) <= d((i + 1) * COL_WIDTH - 1 downto i * COL_WIDTH);
                end if;
            end loop;
        end if;
    end process;

end arch;
